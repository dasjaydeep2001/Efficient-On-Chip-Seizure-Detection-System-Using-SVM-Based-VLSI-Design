
`timescale 1 ns / 1 ns 

module firfilt_tb;

// Function definitions
   function signed [11:0] abs;
   input signed [11:0] arg;
   begin
     abs = arg > 0 ? arg : -arg;
   end
   endfunction // function abs

  task filter_in_data_log_task; 
    input         clk;
    input         reset;
    input         rdenb;
    inout  [9:0]  addr;
    output        done;
  begin

    // Counter to generate the address
    if (reset == 1) 
      addr = 0;
    else begin
      if (rdenb == 1) begin
        if (addr == 999)
          addr = addr; 
        else
          addr =  addr + 1; 
      end
    end

    // Done Signal generation.
    if (reset == 1)
      done = 0; 
    else if (addr == 999)
      done = 1; 
    else
      done = 0; 

  end
  endtask // filter_in_data_log_task

  task filter_out_task; 
    input         clk;
    input         reset;
    input         rdenb;
    inout  [9:0]  addr;
    output        done;
  begin

    // Counter to generate the address
    if (reset == 1) 
      addr = 0;
    else begin
      if (rdenb == 1) begin
        if (addr == 999)
          addr = addr; 
        else
          addr = #1  addr + 1; 
      end
    end

    // Done Signal generation.
    if (reset == 1)
      done = 0; 
    else if (addr == 999)
      done = 1; 
    else
      done = 0; 

  end
  endtask // filter_out_task

 // Constants
 parameter clk_high                         = 5;
 parameter clk_low                          = 5;
 parameter clk_period                       = 10;
 parameter clk_hold                         = 2;
// -------------------------------------------------------------
//
// Module: firfilt_tb_data
// Generated by MATLAB(R) 9.2 and the Filter Design HDL Coder 3.1.1.
// Generated on: 2018-11-01 17:25:28
// -------------------------------------------------------------

 reg  signed [15:0] filter_in_data_log_force [0:999];
 reg  signed [11:0] filter_out_expected [0:999];


// **************************************
 initial //Input & Output data
 begin

 // Input data for filter_in_data_log
 filter_in_data_log_force[  0] <= 16'h8000;
 filter_in_data_log_force[  1] <= 16'h8000;
 filter_in_data_log_force[  2] <= 16'h7fff;
 filter_in_data_log_force[  3] <= 16'h7fff;
 filter_in_data_log_force[  4] <= 16'h8000;
 filter_in_data_log_force[  5] <= 16'h8000;
 filter_in_data_log_force[  6] <= 16'h7fff;
 filter_in_data_log_force[  7] <= 16'h8000;
 filter_in_data_log_force[  8] <= 16'h8000;
 filter_in_data_log_force[  9] <= 16'h7fff;
 filter_in_data_log_force[ 10] <= 16'h8000;
 filter_in_data_log_force[ 11] <= 16'h8000;
 filter_in_data_log_force[ 12] <= 16'h7fff;
 filter_in_data_log_force[ 13] <= 16'h8000;
 filter_in_data_log_force[ 14] <= 16'h8000;
 filter_in_data_log_force[ 15] <= 16'h7fff;
 filter_in_data_log_force[ 16] <= 16'h7fff;
 filter_in_data_log_force[ 17] <= 16'h8000;
 filter_in_data_log_force[ 18] <= 16'h8000;
 filter_in_data_log_force[ 19] <= 16'h7fff;
 filter_in_data_log_force[ 20] <= 16'h8000;
 filter_in_data_log_force[ 21] <= 16'h8000;
 filter_in_data_log_force[ 22] <= 16'h7fff;
 filter_in_data_log_force[ 23] <= 16'h8000;
 filter_in_data_log_force[ 24] <= 16'h8000;
 filter_in_data_log_force[ 25] <= 16'h7fff;
 filter_in_data_log_force[ 26] <= 16'h7fff;
 filter_in_data_log_force[ 27] <= 16'h8000;
 filter_in_data_log_force[ 28] <= 16'h7fff;
 filter_in_data_log_force[ 29] <= 16'h7fff;
 filter_in_data_log_force[ 30] <= 16'h8000;
 filter_in_data_log_force[ 31] <= 16'h8000;
 filter_in_data_log_force[ 32] <= 16'h7fff;
 filter_in_data_log_force[ 33] <= 16'h8000;
 filter_in_data_log_force[ 34] <= 16'h8000;
 filter_in_data_log_force[ 35] <= 16'h8000;
 filter_in_data_log_force[ 36] <= 16'h8000;
 filter_in_data_log_force[ 37] <= 16'h7fff;
 filter_in_data_log_force[ 38] <= 16'h7fff;
 filter_in_data_log_force[ 39] <= 16'h7fff;
 filter_in_data_log_force[ 40] <= 16'h8000;
 filter_in_data_log_force[ 41] <= 16'h8000;
 filter_in_data_log_force[ 42] <= 16'h8000;
 filter_in_data_log_force[ 43] <= 16'h8000;
 filter_in_data_log_force[ 44] <= 16'h8000;
 filter_in_data_log_force[ 45] <= 16'h7fff;
 filter_in_data_log_force[ 46] <= 16'h8000;
 filter_in_data_log_force[ 47] <= 16'h8000;
 filter_in_data_log_force[ 48] <= 16'h7fff;
 filter_in_data_log_force[ 49] <= 16'h8000;
 filter_in_data_log_force[ 50] <= 16'h8000;
 filter_in_data_log_force[ 51] <= 16'h7fff;
 filter_in_data_log_force[ 52] <= 16'h7fff;
 filter_in_data_log_force[ 53] <= 16'h8000;
 filter_in_data_log_force[ 54] <= 16'h8000;
 filter_in_data_log_force[ 55] <= 16'h7fff;
 filter_in_data_log_force[ 56] <= 16'h8000;
 filter_in_data_log_force[ 57] <= 16'h8000;
 filter_in_data_log_force[ 58] <= 16'h7fff;
 filter_in_data_log_force[ 59] <= 16'h7fff;
 filter_in_data_log_force[ 60] <= 16'h8000;
 filter_in_data_log_force[ 61] <= 16'h7fff;
 filter_in_data_log_force[ 62] <= 16'h7fff;
 filter_in_data_log_force[ 63] <= 16'h8000;
 filter_in_data_log_force[ 64] <= 16'h7fff;
 filter_in_data_log_force[ 65] <= 16'h7fff;
 filter_in_data_log_force[ 66] <= 16'h7fff;
 filter_in_data_log_force[ 67] <= 16'h7fff;
 filter_in_data_log_force[ 68] <= 16'h7fff;
 filter_in_data_log_force[ 69] <= 16'h7fff;
 filter_in_data_log_force[ 70] <= 16'h8000;
 filter_in_data_log_force[ 71] <= 16'h7fff;
 filter_in_data_log_force[ 72] <= 16'h7fff;
 filter_in_data_log_force[ 73] <= 16'h8000;
 filter_in_data_log_force[ 74] <= 16'h7fff;
 filter_in_data_log_force[ 75] <= 16'h7fff;
 filter_in_data_log_force[ 76] <= 16'h8000;
 filter_in_data_log_force[ 77] <= 16'h7fff;
 filter_in_data_log_force[ 78] <= 16'h7fff;
 filter_in_data_log_force[ 79] <= 16'h8000;
 filter_in_data_log_force[ 80] <= 16'h8000;
 filter_in_data_log_force[ 81] <= 16'h7fff;
 filter_in_data_log_force[ 82] <= 16'h8000;
 filter_in_data_log_force[ 83] <= 16'h8000;
 filter_in_data_log_force[ 84] <= 16'h7fff;
 filter_in_data_log_force[ 85] <= 16'h7fff;
 filter_in_data_log_force[ 86] <= 16'h8000;
 filter_in_data_log_force[ 87] <= 16'h7fff;
 filter_in_data_log_force[ 88] <= 16'h7fff;
 filter_in_data_log_force[ 89] <= 16'h8000;
 filter_in_data_log_force[ 90] <= 16'h8000;
 filter_in_data_log_force[ 91] <= 16'h7fff;
 filter_in_data_log_force[ 92] <= 16'h8000;
 filter_in_data_log_force[ 93] <= 16'h8000;
 filter_in_data_log_force[ 94] <= 16'h7fff;
 filter_in_data_log_force[ 95] <= 16'h8000;
 filter_in_data_log_force[ 96] <= 16'h8000;
 filter_in_data_log_force[ 97] <= 16'h7fff;
 filter_in_data_log_force[ 98] <= 16'h7fff;
 filter_in_data_log_force[ 99] <= 16'h8000;
 filter_in_data_log_force[100] <= 16'h7fff;
 filter_in_data_log_force[101] <= 16'h7fff;
 filter_in_data_log_force[102] <= 16'h8000;
 filter_in_data_log_force[103] <= 16'h8000;
 filter_in_data_log_force[104] <= 16'h7fff;
 filter_in_data_log_force[105] <= 16'h8000;
 filter_in_data_log_force[106] <= 16'h8000;
 filter_in_data_log_force[107] <= 16'h7fff;
 filter_in_data_log_force[108] <= 16'h8000;
 filter_in_data_log_force[109] <= 16'h8000;
 filter_in_data_log_force[110] <= 16'h7fff;
 filter_in_data_log_force[111] <= 16'h7fff;
 filter_in_data_log_force[112] <= 16'h8000;
 filter_in_data_log_force[113] <= 16'h7fff;
 filter_in_data_log_force[114] <= 16'h7fff;
 filter_in_data_log_force[115] <= 16'h8000;
 filter_in_data_log_force[116] <= 16'h8000;
 filter_in_data_log_force[117] <= 16'h7fff;
 filter_in_data_log_force[118] <= 16'h8000;
 filter_in_data_log_force[119] <= 16'h8000;
 filter_in_data_log_force[120] <= 16'h7fff;
 filter_in_data_log_force[121] <= 16'h8000;
 filter_in_data_log_force[122] <= 16'h8000;
 filter_in_data_log_force[123] <= 16'h8000;
 filter_in_data_log_force[124] <= 16'h8000;
 filter_in_data_log_force[125] <= 16'h8000;
 filter_in_data_log_force[126] <= 16'h7fff;
 filter_in_data_log_force[127] <= 16'h7fff;
 filter_in_data_log_force[128] <= 16'h7fff;
 filter_in_data_log_force[129] <= 16'h8000;
 filter_in_data_log_force[130] <= 16'h8000;
 filter_in_data_log_force[131] <= 16'h8000;
 filter_in_data_log_force[132] <= 16'h8000;
 filter_in_data_log_force[133] <= 16'h7fff;
 filter_in_data_log_force[134] <= 16'h8000;
 filter_in_data_log_force[135] <= 16'h8000;
 filter_in_data_log_force[136] <= 16'h8000;
 filter_in_data_log_force[137] <= 16'h7fff;
 filter_in_data_log_force[138] <= 16'h8000;
 filter_in_data_log_force[139] <= 16'h8000;
 filter_in_data_log_force[140] <= 16'h7fff;
 filter_in_data_log_force[141] <= 16'h8000;
 filter_in_data_log_force[142] <= 16'h8000;
 filter_in_data_log_force[143] <= 16'h7fff;
 filter_in_data_log_force[144] <= 16'h7fff;
 filter_in_data_log_force[145] <= 16'h8000;
 filter_in_data_log_force[146] <= 16'h7fff;
 filter_in_data_log_force[147] <= 16'h7fff;
 filter_in_data_log_force[148] <= 16'h8000;
 filter_in_data_log_force[149] <= 16'h7fff;
 filter_in_data_log_force[150] <= 16'h7fff;
 filter_in_data_log_force[151] <= 16'h7fff;
 filter_in_data_log_force[152] <= 16'h7fff;
 filter_in_data_log_force[153] <= 16'h7fff;
 filter_in_data_log_force[154] <= 16'h7fff;
 filter_in_data_log_force[155] <= 16'h7fff;
 filter_in_data_log_force[156] <= 16'h7fff;
 filter_in_data_log_force[157] <= 16'h7fff;
 filter_in_data_log_force[158] <= 16'h8000;
 filter_in_data_log_force[159] <= 16'h7fff;
 filter_in_data_log_force[160] <= 16'h7fff;
 filter_in_data_log_force[161] <= 16'h8000;
 filter_in_data_log_force[162] <= 16'h8000;
 filter_in_data_log_force[163] <= 16'h7fff;
 filter_in_data_log_force[164] <= 16'h8000;
 filter_in_data_log_force[165] <= 16'h8000;
 filter_in_data_log_force[166] <= 16'h7fff;
 filter_in_data_log_force[167] <= 16'h8000;
 filter_in_data_log_force[168] <= 16'h8000;
 filter_in_data_log_force[169] <= 16'h7fff;
 filter_in_data_log_force[170] <= 16'h7fff;
 filter_in_data_log_force[171] <= 16'h8000;
 filter_in_data_log_force[172] <= 16'h7fff;
 filter_in_data_log_force[173] <= 16'h7fff;
 filter_in_data_log_force[174] <= 16'h8000;
 filter_in_data_log_force[175] <= 16'h8000;
 filter_in_data_log_force[176] <= 16'h7fff;
 filter_in_data_log_force[177] <= 16'h8000;
 filter_in_data_log_force[178] <= 16'h8000;
 filter_in_data_log_force[179] <= 16'h7fff;
 filter_in_data_log_force[180] <= 16'h8000;
 filter_in_data_log_force[181] <= 16'h8000;
 filter_in_data_log_force[182] <= 16'h7fff;
 filter_in_data_log_force[183] <= 16'h7fff;
 filter_in_data_log_force[184] <= 16'h8000;
 filter_in_data_log_force[185] <= 16'h8000;
 filter_in_data_log_force[186] <= 16'h7fff;
 filter_in_data_log_force[187] <= 16'h8000;
 filter_in_data_log_force[188] <= 16'h8000;
 filter_in_data_log_force[189] <= 16'h7fff;
 filter_in_data_log_force[190] <= 16'h8000;
 filter_in_data_log_force[191] <= 16'h8000;
 filter_in_data_log_force[192] <= 16'h7fff;
 filter_in_data_log_force[193] <= 16'h8000;
 filter_in_data_log_force[194] <= 16'h8000;
 filter_in_data_log_force[195] <= 16'h7fff;
 filter_in_data_log_force[196] <= 16'h7fff;
 filter_in_data_log_force[197] <= 16'h8000;
 filter_in_data_log_force[198] <= 16'h7fff;
 filter_in_data_log_force[199] <= 16'h7fff;
 filter_in_data_log_force[200] <= 16'h8000;
 filter_in_data_log_force[201] <= 16'h8000;
 filter_in_data_log_force[202] <= 16'h7fff;
 filter_in_data_log_force[203] <= 16'h8000;
 filter_in_data_log_force[204] <= 16'h8000;
 filter_in_data_log_force[205] <= 16'h7fff;
 filter_in_data_log_force[206] <= 16'h8000;
 filter_in_data_log_force[207] <= 16'h8000;
 filter_in_data_log_force[208] <= 16'h8000;
 filter_in_data_log_force[209] <= 16'h7fff;
 filter_in_data_log_force[210] <= 16'h7fff;
 filter_in_data_log_force[211] <= 16'h7fff;
 filter_in_data_log_force[212] <= 16'h7fff;
 filter_in_data_log_force[213] <= 16'h8000;
 filter_in_data_log_force[214] <= 16'h8000;
 filter_in_data_log_force[215] <= 16'h8000;
 filter_in_data_log_force[216] <= 16'h8000;
 filter_in_data_log_force[217] <= 16'h8000;
 filter_in_data_log_force[218] <= 16'h7fff;
 filter_in_data_log_force[219] <= 16'h8000;
 filter_in_data_log_force[220] <= 16'h8000;
 filter_in_data_log_force[221] <= 16'h8000;
 filter_in_data_log_force[222] <= 16'h7fff;
 filter_in_data_log_force[223] <= 16'h8000;
 filter_in_data_log_force[224] <= 16'h8000;
 filter_in_data_log_force[225] <= 16'h7fff;
 filter_in_data_log_force[226] <= 16'h8000;
 filter_in_data_log_force[227] <= 16'h8000;
 filter_in_data_log_force[228] <= 16'h7fff;
 filter_in_data_log_force[229] <= 16'h7fff;
 filter_in_data_log_force[230] <= 16'h8000;
 filter_in_data_log_force[231] <= 16'h7fff;
 filter_in_data_log_force[232] <= 16'h7fff;
 filter_in_data_log_force[233] <= 16'h8000;
 filter_in_data_log_force[234] <= 16'h7fff;
 filter_in_data_log_force[235] <= 16'h7fff;
 filter_in_data_log_force[236] <= 16'h7fff;
 filter_in_data_log_force[237] <= 16'h7fff;
 filter_in_data_log_force[238] <= 16'h7fff;
 filter_in_data_log_force[239] <= 16'h7fff;
 filter_in_data_log_force[240] <= 16'hd970;
 filter_in_data_log_force[241] <= 16'h7fff;
 filter_in_data_log_force[242] <= 16'h7fff;
 filter_in_data_log_force[243] <= 16'h8000;
 filter_in_data_log_force[244] <= 16'h7fff;
 filter_in_data_log_force[245] <= 16'h7fff;
 filter_in_data_log_force[246] <= 16'h8000;
 filter_in_data_log_force[247] <= 16'h8000;
 filter_in_data_log_force[248] <= 16'h7fff;
 filter_in_data_log_force[249] <= 16'h8000;
 filter_in_data_log_force[250] <= 16'h8000;
 filter_in_data_log_force[251] <= 16'h7fff;
 filter_in_data_log_force[252] <= 16'h8000;
 filter_in_data_log_force[253] <= 16'h8000;
 filter_in_data_log_force[254] <= 16'h7fff;
 filter_in_data_log_force[255] <= 16'h7fff;
 filter_in_data_log_force[256] <= 16'h8000;
 filter_in_data_log_force[257] <= 16'h5759;
 filter_in_data_log_force[258] <= 16'h7fff;
 filter_in_data_log_force[259] <= 16'h8000;
 filter_in_data_log_force[260] <= 16'h8000;
 filter_in_data_log_force[261] <= 16'h7fff;
 filter_in_data_log_force[262] <= 16'h8000;
 filter_in_data_log_force[263] <= 16'h8000;
 filter_in_data_log_force[264] <= 16'h7fff;
 filter_in_data_log_force[265] <= 16'h8000;
 filter_in_data_log_force[266] <= 16'h8000;
 filter_in_data_log_force[267] <= 16'h7fff;
 filter_in_data_log_force[268] <= 16'h7fff;
 filter_in_data_log_force[269] <= 16'h8000;
 filter_in_data_log_force[270] <= 16'h8000;
 filter_in_data_log_force[271] <= 16'h7fff;
 filter_in_data_log_force[272] <= 16'h8000;
 filter_in_data_log_force[273] <= 16'h8000;
 filter_in_data_log_force[274] <= 16'h7fff;
 filter_in_data_log_force[275] <= 16'h8000;
 filter_in_data_log_force[276] <= 16'h8000;
 filter_in_data_log_force[277] <= 16'h7fff;
 filter_in_data_log_force[278] <= 16'h7fff;
 filter_in_data_log_force[279] <= 16'h8000;
 filter_in_data_log_force[280] <= 16'h7fff;
 filter_in_data_log_force[281] <= 16'h7fff;
 filter_in_data_log_force[282] <= 16'h8000;
 filter_in_data_log_force[283] <= 16'h28a7;
 filter_in_data_log_force[284] <= 16'h7fff;
 filter_in_data_log_force[285] <= 16'h8000;
 filter_in_data_log_force[286] <= 16'h8000;
 filter_in_data_log_force[287] <= 16'h7fff;
 filter_in_data_log_force[288] <= 16'h8000;
 filter_in_data_log_force[289] <= 16'h8000;
 filter_in_data_log_force[290] <= 16'h8000;
 filter_in_data_log_force[291] <= 16'h8000;
 filter_in_data_log_force[292] <= 16'h8000;
 filter_in_data_log_force[293] <= 16'h7fff;
 filter_in_data_log_force[294] <= 16'h7fff;
 filter_in_data_log_force[295] <= 16'h7fff;
 filter_in_data_log_force[296] <= 16'h8000;
 filter_in_data_log_force[297] <= 16'h8000;
 filter_in_data_log_force[298] <= 16'h8000;
 filter_in_data_log_force[299] <= 16'h8000;
 filter_in_data_log_force[300] <= 16'h7fff;
 filter_in_data_log_force[301] <= 16'h8000;
 filter_in_data_log_force[302] <= 16'h8000;
 filter_in_data_log_force[303] <= 16'h8000;
 filter_in_data_log_force[304] <= 16'h7fff;
 filter_in_data_log_force[305] <= 16'h8000;
 filter_in_data_log_force[306] <= 16'h8000;
 filter_in_data_log_force[307] <= 16'h7fff;
 filter_in_data_log_force[308] <= 16'h8000;
 filter_in_data_log_force[309] <= 16'h8000;
 filter_in_data_log_force[310] <= 16'h7fff;
 filter_in_data_log_force[311] <= 16'h8000;
 filter_in_data_log_force[312] <= 16'h8000;
 filter_in_data_log_force[313] <= 16'h7fff;
 filter_in_data_log_force[314] <= 16'h7fff;
 filter_in_data_log_force[315] <= 16'h8000;
 filter_in_data_log_force[316] <= 16'h7fff;
 filter_in_data_log_force[317] <= 16'h7fff;
 filter_in_data_log_force[318] <= 16'h7fff;
 filter_in_data_log_force[319] <= 16'h7fff;
 filter_in_data_log_force[320] <= 16'h7fff;
 filter_in_data_log_force[321] <= 16'h7fff;
 filter_in_data_log_force[322] <= 16'h7fff;
 filter_in_data_log_force[323] <= 16'h7fff;
 filter_in_data_log_force[324] <= 16'h7fff;
 filter_in_data_log_force[325] <= 16'h8000;
 filter_in_data_log_force[326] <= 16'h7fff;
 filter_in_data_log_force[327] <= 16'h7fff;
 filter_in_data_log_force[328] <= 16'h8000;
 filter_in_data_log_force[329] <= 16'h7fff;
 filter_in_data_log_force[330] <= 16'h7fff;
 filter_in_data_log_force[331] <= 16'h8000;
 filter_in_data_log_force[332] <= 16'h8000;
 filter_in_data_log_force[333] <= 16'h7fff;
 filter_in_data_log_force[334] <= 16'h8000;
 filter_in_data_log_force[335] <= 16'h8000;
 filter_in_data_log_force[336] <= 16'h7fff;
 filter_in_data_log_force[337] <= 16'h5759;
 filter_in_data_log_force[338] <= 16'h8000;
 filter_in_data_log_force[339] <= 16'h7fff;
 filter_in_data_log_force[340] <= 16'h7fff;
 filter_in_data_log_force[341] <= 16'h8000;
 filter_in_data_log_force[342] <= 16'h8000;
 filter_in_data_log_force[343] <= 16'h7fff;
 filter_in_data_log_force[344] <= 16'h8000;
 filter_in_data_log_force[345] <= 16'h8000;
 filter_in_data_log_force[346] <= 16'h7fff;
 filter_in_data_log_force[347] <= 16'h8000;
 filter_in_data_log_force[348] <= 16'h8000;
 filter_in_data_log_force[349] <= 16'h7fff;
 filter_in_data_log_force[350] <= 16'h8000;
 filter_in_data_log_force[351] <= 16'h8000;
 filter_in_data_log_force[352] <= 16'h8000;
 filter_in_data_log_force[353] <= 16'h7fff;
 filter_in_data_log_force[354] <= 16'h8000;
 filter_in_data_log_force[355] <= 16'h8000;
 filter_in_data_log_force[356] <= 16'h7fff;
 filter_in_data_log_force[357] <= 16'h8000;
 filter_in_data_log_force[358] <= 16'h8000;
 filter_in_data_log_force[359] <= 16'h7fff;
 filter_in_data_log_force[360] <= 16'h8000;
 filter_in_data_log_force[361] <= 16'h8000;
 filter_in_data_log_force[362] <= 16'h7fff;
 filter_in_data_log_force[363] <= 16'h7fff;
 filter_in_data_log_force[364] <= 16'h8000;
 filter_in_data_log_force[365] <= 16'h7fff;
 filter_in_data_log_force[366] <= 16'h7fff;
 filter_in_data_log_force[367] <= 16'h8000;
 filter_in_data_log_force[368] <= 16'h8000;
 filter_in_data_log_force[369] <= 16'h7fff;
 filter_in_data_log_force[370] <= 16'h8000;
 filter_in_data_log_force[371] <= 16'h8000;
 filter_in_data_log_force[372] <= 16'h7fff;
 filter_in_data_log_force[373] <= 16'h8000;
 filter_in_data_log_force[374] <= 16'h8000;
 filter_in_data_log_force[375] <= 16'h7fff;
 filter_in_data_log_force[376] <= 16'h7fff;
 filter_in_data_log_force[377] <= 16'h7fff;
 filter_in_data_log_force[378] <= 16'h7fff;
 filter_in_data_log_force[379] <= 16'h8000;
 filter_in_data_log_force[380] <= 16'h8000;
 filter_in_data_log_force[381] <= 16'h8000;
 filter_in_data_log_force[382] <= 16'h7fff;
 filter_in_data_log_force[383] <= 16'h8000;
 filter_in_data_log_force[384] <= 16'h8000;
 filter_in_data_log_force[385] <= 16'h7fff;
 filter_in_data_log_force[386] <= 16'h8000;
 filter_in_data_log_force[387] <= 16'h8000;
 filter_in_data_log_force[388] <= 16'h8000;
 filter_in_data_log_force[389] <= 16'h7fff;
 filter_in_data_log_force[390] <= 16'h8000;
 filter_in_data_log_force[391] <= 16'h8000;
 filter_in_data_log_force[392] <= 16'h7fff;
 filter_in_data_log_force[393] <= 16'h8000;
 filter_in_data_log_force[394] <= 16'h8000;
 filter_in_data_log_force[395] <= 16'h7fff;
 filter_in_data_log_force[396] <= 16'h7fff;
 filter_in_data_log_force[397] <= 16'h8000;
 filter_in_data_log_force[398] <= 16'h7fff;
 filter_in_data_log_force[399] <= 16'h7fff;
 filter_in_data_log_force[400] <= 16'h8000;
 filter_in_data_log_force[401] <= 16'h7fff;
 filter_in_data_log_force[402] <= 16'h7fff;
 filter_in_data_log_force[403] <= 16'h7fff;
 filter_in_data_log_force[404] <= 16'h7fff;
 filter_in_data_log_force[405] <= 16'h7fff;
 filter_in_data_log_force[406] <= 16'h7fff;
 filter_in_data_log_force[407] <= 16'h8000;
 filter_in_data_log_force[408] <= 16'h7fff;
 filter_in_data_log_force[409] <= 16'h7fff;
 filter_in_data_log_force[410] <= 16'h8000;
 filter_in_data_log_force[411] <= 16'h7fff;
 filter_in_data_log_force[412] <= 16'h7fff;
 filter_in_data_log_force[413] <= 16'h8000;
 filter_in_data_log_force[414] <= 16'h8000;
 filter_in_data_log_force[415] <= 16'h7fff;
 filter_in_data_log_force[416] <= 16'h8000;
 filter_in_data_log_force[417] <= 16'h8000;
 filter_in_data_log_force[418] <= 16'h7fff;
 filter_in_data_log_force[419] <= 16'h8000;
 filter_in_data_log_force[420] <= 16'h8000;
 filter_in_data_log_force[421] <= 16'h7fff;
 filter_in_data_log_force[422] <= 16'h7fff;
 filter_in_data_log_force[423] <= 16'h8000;
 filter_in_data_log_force[424] <= 16'h7fff;
 filter_in_data_log_force[425] <= 16'h7fff;
 filter_in_data_log_force[426] <= 16'h8000;
 filter_in_data_log_force[427] <= 16'h8000;
 filter_in_data_log_force[428] <= 16'h7fff;
 filter_in_data_log_force[429] <= 16'h8000;
 filter_in_data_log_force[430] <= 16'h8000;
 filter_in_data_log_force[431] <= 16'h7fff;
 filter_in_data_log_force[432] <= 16'h8000;
 filter_in_data_log_force[433] <= 16'h8000;
 filter_in_data_log_force[434] <= 16'h7fff;
 filter_in_data_log_force[435] <= 16'h7fff;
 filter_in_data_log_force[436] <= 16'h8000;
 filter_in_data_log_force[437] <= 16'h8000;
 filter_in_data_log_force[438] <= 16'h7fff;
 filter_in_data_log_force[439] <= 16'h8000;
 filter_in_data_log_force[440] <= 16'h8000;
 filter_in_data_log_force[441] <= 16'h7fff;
 filter_in_data_log_force[442] <= 16'h8000;
 filter_in_data_log_force[443] <= 16'h8000;
 filter_in_data_log_force[444] <= 16'h7fff;
 filter_in_data_log_force[445] <= 16'h8000;
 filter_in_data_log_force[446] <= 16'h8000;
 filter_in_data_log_force[447] <= 16'h7fff;
 filter_in_data_log_force[448] <= 16'h7fff;
 filter_in_data_log_force[449] <= 16'h8000;
 filter_in_data_log_force[450] <= 16'h7fff;
 filter_in_data_log_force[451] <= 16'h7fff;
 filter_in_data_log_force[452] <= 16'h8000;
 filter_in_data_log_force[453] <= 16'h8000;
 filter_in_data_log_force[454] <= 16'h7fff;
 filter_in_data_log_force[455] <= 16'h8000;
 filter_in_data_log_force[456] <= 16'h8000;
 filter_in_data_log_force[457] <= 16'h7fff;
 filter_in_data_log_force[458] <= 16'h8000;
 filter_in_data_log_force[459] <= 16'h8000;
 filter_in_data_log_force[460] <= 16'h8000;
 filter_in_data_log_force[461] <= 16'h8000;
 filter_in_data_log_force[462] <= 16'h8000;
 filter_in_data_log_force[463] <= 16'h7fff;
 filter_in_data_log_force[464] <= 16'h7fff;
 filter_in_data_log_force[465] <= 16'h7fff;
 filter_in_data_log_force[466] <= 16'h8000;
 filter_in_data_log_force[467] <= 16'h8000;
 filter_in_data_log_force[468] <= 16'h8000;
 filter_in_data_log_force[469] <= 16'h8000;
 filter_in_data_log_force[470] <= 16'h7fff;
 filter_in_data_log_force[471] <= 16'h8000;
 filter_in_data_log_force[472] <= 16'h8000;
 filter_in_data_log_force[473] <= 16'h8000;
 filter_in_data_log_force[474] <= 16'h7fff;
 filter_in_data_log_force[475] <= 16'h8000;
 filter_in_data_log_force[476] <= 16'h8000;
 filter_in_data_log_force[477] <= 16'h7fff;
 filter_in_data_log_force[478] <= 16'h8000;
 filter_in_data_log_force[479] <= 16'h8000;
 filter_in_data_log_force[480] <= 16'h7fff;
 filter_in_data_log_force[481] <= 16'h7fff;
 filter_in_data_log_force[482] <= 16'h8000;
 filter_in_data_log_force[483] <= 16'h7fff;
 filter_in_data_log_force[484] <= 16'h7fff;
 filter_in_data_log_force[485] <= 16'h8000;
 filter_in_data_log_force[486] <= 16'h7fff;
 filter_in_data_log_force[487] <= 16'h7fff;
 filter_in_data_log_force[488] <= 16'h7fff;
 filter_in_data_log_force[489] <= 16'h7fff;
 filter_in_data_log_force[490] <= 16'h7fff;
 filter_in_data_log_force[491] <= 16'h7fff;
 filter_in_data_log_force[492] <= 16'h7fff;
 filter_in_data_log_force[493] <= 16'h7fff;
 filter_in_data_log_force[494] <= 16'h7fff;
 filter_in_data_log_force[495] <= 16'h8000;
 filter_in_data_log_force[496] <= 16'h7fff;
 filter_in_data_log_force[497] <= 16'h7fff;
 filter_in_data_log_force[498] <= 16'h8000;
 filter_in_data_log_force[499] <= 16'h8000;
 filter_in_data_log_force[500] <= 16'h7fff;
 filter_in_data_log_force[501] <= 16'h8000;
 filter_in_data_log_force[502] <= 16'h8000;
 filter_in_data_log_force[503] <= 16'h7fff;
 filter_in_data_log_force[504] <= 16'h7fff;
 filter_in_data_log_force[505] <= 16'h8000;
 filter_in_data_log_force[506] <= 16'h7fff;
 filter_in_data_log_force[507] <= 16'h7fff;
 filter_in_data_log_force[508] <= 16'h8000;
 filter_in_data_log_force[509] <= 16'h7fff;
 filter_in_data_log_force[510] <= 16'h7fff;
 filter_in_data_log_force[511] <= 16'h8000;
 filter_in_data_log_force[512] <= 16'h8000;
 filter_in_data_log_force[513] <= 16'h7fff;
 filter_in_data_log_force[514] <= 16'h8000;
 filter_in_data_log_force[515] <= 16'h8000;
 filter_in_data_log_force[516] <= 16'h7fff;
 filter_in_data_log_force[517] <= 16'h7fff;
 filter_in_data_log_force[518] <= 16'h8000;
 filter_in_data_log_force[519] <= 16'h7fff;
 filter_in_data_log_force[520] <= 16'h7fff;
 filter_in_data_log_force[521] <= 16'h8000;
 filter_in_data_log_force[522] <= 16'h8000;
 filter_in_data_log_force[523] <= 16'h7fff;
 filter_in_data_log_force[524] <= 16'h8000;
 filter_in_data_log_force[525] <= 16'h8000;
 filter_in_data_log_force[526] <= 16'h7fff;
 filter_in_data_log_force[527] <= 16'h8000;
 filter_in_data_log_force[528] <= 16'h8000;
 filter_in_data_log_force[529] <= 16'h7fff;
 filter_in_data_log_force[530] <= 16'h7fff;
 filter_in_data_log_force[531] <= 16'h8000;
 filter_in_data_log_force[532] <= 16'h7fff;
 filter_in_data_log_force[533] <= 16'h7fff;
 filter_in_data_log_force[534] <= 16'h8000;
 filter_in_data_log_force[535] <= 16'h8000;
 filter_in_data_log_force[536] <= 16'h7fff;
 filter_in_data_log_force[537] <= 16'h8000;
 filter_in_data_log_force[538] <= 16'h8000;
 filter_in_data_log_force[539] <= 16'h7fff;
 filter_in_data_log_force[540] <= 16'h8000;
 filter_in_data_log_force[541] <= 16'h8000;
 filter_in_data_log_force[542] <= 16'h7fff;
 filter_in_data_log_force[543] <= 16'h7fff;
 filter_in_data_log_force[544] <= 16'h8000;
 filter_in_data_log_force[545] <= 16'h7fff;
 filter_in_data_log_force[546] <= 16'h7fff;
 filter_in_data_log_force[547] <= 16'h8000;
 filter_in_data_log_force[548] <= 16'h8000;
 filter_in_data_log_force[549] <= 16'h7fff;
 filter_in_data_log_force[550] <= 16'h8000;
 filter_in_data_log_force[551] <= 16'h8000;
 filter_in_data_log_force[552] <= 16'h7fff;
 filter_in_data_log_force[553] <= 16'h8000;
 filter_in_data_log_force[554] <= 16'h8000;
 filter_in_data_log_force[555] <= 16'h8000;
 filter_in_data_log_force[556] <= 16'h7fff;
 filter_in_data_log_force[557] <= 16'h7fff;
 filter_in_data_log_force[558] <= 16'h7fff;
 filter_in_data_log_force[559] <= 16'h7fff;
 filter_in_data_log_force[560] <= 16'h8000;
 filter_in_data_log_force[561] <= 16'h8000;
 filter_in_data_log_force[562] <= 16'h8000;
 filter_in_data_log_force[563] <= 16'h8000;
 filter_in_data_log_force[564] <= 16'h8000;
 filter_in_data_log_force[565] <= 16'h7fff;
 filter_in_data_log_force[566] <= 16'h8000;
 filter_in_data_log_force[567] <= 16'h8000;
 filter_in_data_log_force[568] <= 16'h8000;
 filter_in_data_log_force[569] <= 16'h7fff;
 filter_in_data_log_force[570] <= 16'h8000;
 filter_in_data_log_force[571] <= 16'h8000;
 filter_in_data_log_force[572] <= 16'h7fff;
 filter_in_data_log_force[573] <= 16'h8000;
 filter_in_data_log_force[574] <= 16'h8000;
 filter_in_data_log_force[575] <= 16'h7fff;
 filter_in_data_log_force[576] <= 16'h7fff;
 filter_in_data_log_force[577] <= 16'h8000;
 filter_in_data_log_force[578] <= 16'h7fff;
 filter_in_data_log_force[579] <= 16'h7fff;
 filter_in_data_log_force[580] <= 16'h8000;
 filter_in_data_log_force[581] <= 16'h7fff;
 filter_in_data_log_force[582] <= 16'h7fff;
 filter_in_data_log_force[583] <= 16'h7fff;
 filter_in_data_log_force[584] <= 16'h7fff;
 filter_in_data_log_force[585] <= 16'h7fff;
 filter_in_data_log_force[586] <= 16'h7fff;
 filter_in_data_log_force[587] <= 16'h7fff;
 filter_in_data_log_force[588] <= 16'h7fff;
 filter_in_data_log_force[589] <= 16'h7fff;
 filter_in_data_log_force[590] <= 16'h8000;
 filter_in_data_log_force[591] <= 16'h7fff;
 filter_in_data_log_force[592] <= 16'h7fff;
 filter_in_data_log_force[593] <= 16'h8000;
 filter_in_data_log_force[594] <= 16'h7fff;
 filter_in_data_log_force[595] <= 16'h7fff;
 filter_in_data_log_force[596] <= 16'h8000;
 filter_in_data_log_force[597] <= 16'h8000;
 filter_in_data_log_force[598] <= 16'h7fff;
 filter_in_data_log_force[599] <= 16'h8000;
 filter_in_data_log_force[600] <= 16'h8000;
 filter_in_data_log_force[601] <= 16'h7fff;
 filter_in_data_log_force[602] <= 16'h7fff;
 filter_in_data_log_force[603] <= 16'h8000;
 filter_in_data_log_force[604] <= 16'h7fff;
 filter_in_data_log_force[605] <= 16'h7fff;
 filter_in_data_log_force[606] <= 16'h8000;
 filter_in_data_log_force[607] <= 16'h8000;
 filter_in_data_log_force[608] <= 16'h7fff;
 filter_in_data_log_force[609] <= 16'h8000;
 filter_in_data_log_force[610] <= 16'h8000;
 filter_in_data_log_force[611] <= 16'h7fff;
 filter_in_data_log_force[612] <= 16'h8000;
 filter_in_data_log_force[613] <= 16'h8000;
 filter_in_data_log_force[614] <= 16'h7fff;
 filter_in_data_log_force[615] <= 16'h7fff;
 filter_in_data_log_force[616] <= 16'h8000;
 filter_in_data_log_force[617] <= 16'h8000;
 filter_in_data_log_force[618] <= 16'h7fff;
 filter_in_data_log_force[619] <= 16'h8000;
 filter_in_data_log_force[620] <= 16'h8000;
 filter_in_data_log_force[621] <= 16'h7fff;
 filter_in_data_log_force[622] <= 16'h8000;
 filter_in_data_log_force[623] <= 16'h8000;
 filter_in_data_log_force[624] <= 16'h7fff;
 filter_in_data_log_force[625] <= 16'h8000;
 filter_in_data_log_force[626] <= 16'h8000;
 filter_in_data_log_force[627] <= 16'h7fff;
 filter_in_data_log_force[628] <= 16'h7fff;
 filter_in_data_log_force[629] <= 16'h8000;
 filter_in_data_log_force[630] <= 16'h8000;
 filter_in_data_log_force[631] <= 16'h7fff;
 filter_in_data_log_force[632] <= 16'h8000;
 filter_in_data_log_force[633] <= 16'h8000;
 filter_in_data_log_force[634] <= 16'h7fff;
 filter_in_data_log_force[635] <= 16'h8000;
 filter_in_data_log_force[636] <= 16'h8000;
 filter_in_data_log_force[637] <= 16'h7fff;
 filter_in_data_log_force[638] <= 16'h7fff;
 filter_in_data_log_force[639] <= 16'h8000;
 filter_in_data_log_force[640] <= 16'h7fff;
 filter_in_data_log_force[641] <= 16'h7fff;
 filter_in_data_log_force[642] <= 16'h8000;
 filter_in_data_log_force[643] <= 16'h7fff;
 filter_in_data_log_force[644] <= 16'h7fff;
 filter_in_data_log_force[645] <= 16'h8000;
 filter_in_data_log_force[646] <= 16'h8000;
 filter_in_data_log_force[647] <= 16'h7fff;
 filter_in_data_log_force[648] <= 16'h8000;
 filter_in_data_log_force[649] <= 16'h8000;
 filter_in_data_log_force[650] <= 16'h8000;
 filter_in_data_log_force[651] <= 16'h8000;
 filter_in_data_log_force[652] <= 16'h8000;
 filter_in_data_log_force[653] <= 16'h8000;
 filter_in_data_log_force[654] <= 16'h7fff;
 filter_in_data_log_force[655] <= 16'h7fff;
 filter_in_data_log_force[656] <= 16'h7fff;
 filter_in_data_log_force[657] <= 16'h7fff;
 filter_in_data_log_force[658] <= 16'h8000;
 filter_in_data_log_force[659] <= 16'h8000;
 filter_in_data_log_force[660] <= 16'h8000;
 filter_in_data_log_force[661] <= 16'h8000;
 filter_in_data_log_force[662] <= 16'h8000;
 filter_in_data_log_force[663] <= 16'h8000;
 filter_in_data_log_force[664] <= 16'h7fff;
 filter_in_data_log_force[665] <= 16'h8000;
 filter_in_data_log_force[666] <= 16'h8000;
 filter_in_data_log_force[667] <= 16'h7fff;
 filter_in_data_log_force[668] <= 16'h8000;
 filter_in_data_log_force[669] <= 16'h8000;
 filter_in_data_log_force[670] <= 16'h7fff;
 filter_in_data_log_force[671] <= 16'h8000;
 filter_in_data_log_force[672] <= 16'h8000;
 filter_in_data_log_force[673] <= 16'h7fff;
 filter_in_data_log_force[674] <= 16'h7fff;
 filter_in_data_log_force[675] <= 16'h8000;
 filter_in_data_log_force[676] <= 16'h7fff;
 filter_in_data_log_force[677] <= 16'h7fff;
 filter_in_data_log_force[678] <= 16'h8000;
 filter_in_data_log_force[679] <= 16'h7fff;
 filter_in_data_log_force[680] <= 16'h7fff;
 filter_in_data_log_force[681] <= 16'h7fff;
 filter_in_data_log_force[682] <= 16'h7fff;
 filter_in_data_log_force[683] <= 16'h7fff;
 filter_in_data_log_force[684] <= 16'h7fff;
 filter_in_data_log_force[685] <= 16'h8000;
 filter_in_data_log_force[686] <= 16'h7fff;
 filter_in_data_log_force[687] <= 16'h7fff;
 filter_in_data_log_force[688] <= 16'h8000;
 filter_in_data_log_force[689] <= 16'h7fff;
 filter_in_data_log_force[690] <= 16'h7fff;
 filter_in_data_log_force[691] <= 16'h8000;
 filter_in_data_log_force[692] <= 16'h8000;
 filter_in_data_log_force[693] <= 16'h7fff;
 filter_in_data_log_force[694] <= 16'h8000;
 filter_in_data_log_force[695] <= 16'h8000;
 filter_in_data_log_force[696] <= 16'h7fff;
 filter_in_data_log_force[697] <= 16'h7fff;
 filter_in_data_log_force[698] <= 16'h8000;
 filter_in_data_log_force[699] <= 16'h7fff;
 filter_in_data_log_force[700] <= 16'h7fff;
 filter_in_data_log_force[701] <= 16'h8000;
 filter_in_data_log_force[702] <= 16'h8000;
 filter_in_data_log_force[703] <= 16'h7fff;
 filter_in_data_log_force[704] <= 16'h8000;
 filter_in_data_log_force[705] <= 16'h8000;
 filter_in_data_log_force[706] <= 16'h7fff;
 filter_in_data_log_force[707] <= 16'h8000;
 filter_in_data_log_force[708] <= 16'h8000;
 filter_in_data_log_force[709] <= 16'h7fff;
 filter_in_data_log_force[710] <= 16'h7fff;
 filter_in_data_log_force[711] <= 16'h8000;
 filter_in_data_log_force[712] <= 16'h7fff;
 filter_in_data_log_force[713] <= 16'h7fff;
 filter_in_data_log_force[714] <= 16'h8000;
 filter_in_data_log_force[715] <= 16'h8000;
 filter_in_data_log_force[716] <= 16'h7fff;
 filter_in_data_log_force[717] <= 16'h8000;
 filter_in_data_log_force[718] <= 16'h8000;
 filter_in_data_log_force[719] <= 16'h7fff;
 filter_in_data_log_force[720] <= 16'h8000;
 filter_in_data_log_force[721] <= 16'h8000;
 filter_in_data_log_force[722] <= 16'h7fff;
 filter_in_data_log_force[723] <= 16'h7fff;
 filter_in_data_log_force[724] <= 16'h8000;
 filter_in_data_log_force[725] <= 16'h8000;
 filter_in_data_log_force[726] <= 16'h7fff;
 filter_in_data_log_force[727] <= 16'h8000;
 filter_in_data_log_force[728] <= 16'h8000;
 filter_in_data_log_force[729] <= 16'h7fff;
 filter_in_data_log_force[730] <= 16'h8000;
 filter_in_data_log_force[731] <= 16'h8000;
 filter_in_data_log_force[732] <= 16'h7fff;
 filter_in_data_log_force[733] <= 16'h7fff;
 filter_in_data_log_force[734] <= 16'h8000;
 filter_in_data_log_force[735] <= 16'h7fff;
 filter_in_data_log_force[736] <= 16'h7fff;
 filter_in_data_log_force[737] <= 16'h8000;
 filter_in_data_log_force[738] <= 16'h7fff;
 filter_in_data_log_force[739] <= 16'h7fff;
 filter_in_data_log_force[740] <= 16'h8000;
 filter_in_data_log_force[741] <= 16'h8000;
 filter_in_data_log_force[742] <= 16'h7fff;
 filter_in_data_log_force[743] <= 16'h8000;
 filter_in_data_log_force[744] <= 16'h8000;
 filter_in_data_log_force[745] <= 16'h7fff;
 filter_in_data_log_force[746] <= 16'h8000;
 filter_in_data_log_force[747] <= 16'h8000;
 filter_in_data_log_force[748] <= 16'h7fff;
 filter_in_data_log_force[749] <= 16'h7fff;
 filter_in_data_log_force[750] <= 16'h7fff;
 filter_in_data_log_force[751] <= 16'h7fff;
 filter_in_data_log_force[752] <= 16'h8000;
 filter_in_data_log_force[753] <= 16'h8000;
 filter_in_data_log_force[754] <= 16'h8000;
 filter_in_data_log_force[755] <= 16'h7fff;
 filter_in_data_log_force[756] <= 16'h8000;
 filter_in_data_log_force[757] <= 16'h8000;
 filter_in_data_log_force[758] <= 16'h7fff;
 filter_in_data_log_force[759] <= 16'h7fff;
 filter_in_data_log_force[760] <= 16'h8000;
 filter_in_data_log_force[761] <= 16'h8000;
 filter_in_data_log_force[762] <= 16'h7fff;
 filter_in_data_log_force[763] <= 16'h8000;
 filter_in_data_log_force[764] <= 16'h8000;
 filter_in_data_log_force[765] <= 16'h7fff;
 filter_in_data_log_force[766] <= 16'h8000;
 filter_in_data_log_force[767] <= 16'h8000;
 filter_in_data_log_force[768] <= 16'h7fff;
 filter_in_data_log_force[769] <= 16'h7fff;
 filter_in_data_log_force[770] <= 16'h8000;
 filter_in_data_log_force[771] <= 16'h7fff;
 filter_in_data_log_force[772] <= 16'h7fff;
 filter_in_data_log_force[773] <= 16'h8000;
 filter_in_data_log_force[774] <= 16'h7fff;
 filter_in_data_log_force[775] <= 16'h7fff;
 filter_in_data_log_force[776] <= 16'h7fff;
 filter_in_data_log_force[777] <= 16'h7fff;
 filter_in_data_log_force[778] <= 16'h7fff;
 filter_in_data_log_force[779] <= 16'h7fff;
 filter_in_data_log_force[780] <= 16'h8000;
 filter_in_data_log_force[781] <= 16'h7fff;
 filter_in_data_log_force[782] <= 16'h7fff;
 filter_in_data_log_force[783] <= 16'h8000;
 filter_in_data_log_force[784] <= 16'h7fff;
 filter_in_data_log_force[785] <= 16'h7fff;
 filter_in_data_log_force[786] <= 16'h8000;
 filter_in_data_log_force[787] <= 16'h8000;
 filter_in_data_log_force[788] <= 16'h7fff;
 filter_in_data_log_force[789] <= 16'h8000;
 filter_in_data_log_force[790] <= 16'h8000;
 filter_in_data_log_force[791] <= 16'h7fff;
 filter_in_data_log_force[792] <= 16'h8000;
 filter_in_data_log_force[793] <= 16'h8000;
 filter_in_data_log_force[794] <= 16'h7fff;
 filter_in_data_log_force[795] <= 16'h7fff;
 filter_in_data_log_force[796] <= 16'h8000;
 filter_in_data_log_force[797] <= 16'h5759;
 filter_in_data_log_force[798] <= 16'h7fff;
 filter_in_data_log_force[799] <= 16'h8000;
 filter_in_data_log_force[800] <= 16'h8000;
 filter_in_data_log_force[801] <= 16'h7fff;
 filter_in_data_log_force[802] <= 16'h8000;
 filter_in_data_log_force[803] <= 16'h8000;
 filter_in_data_log_force[804] <= 16'h7fff;
 filter_in_data_log_force[805] <= 16'h8000;
 filter_in_data_log_force[806] <= 16'h8000;
 filter_in_data_log_force[807] <= 16'h7fff;
 filter_in_data_log_force[808] <= 16'h7fff;
 filter_in_data_log_force[809] <= 16'h8000;
 filter_in_data_log_force[810] <= 16'h8000;
 filter_in_data_log_force[811] <= 16'h7fff;
 filter_in_data_log_force[812] <= 16'h8000;
 filter_in_data_log_force[813] <= 16'h8000;
 filter_in_data_log_force[814] <= 16'h7fff;
 filter_in_data_log_force[815] <= 16'h8000;
 filter_in_data_log_force[816] <= 16'h8000;
 filter_in_data_log_force[817] <= 16'h7fff;
 filter_in_data_log_force[818] <= 16'h7fff;
 filter_in_data_log_force[819] <= 16'h8000;
 filter_in_data_log_force[820] <= 16'h7fff;
 filter_in_data_log_force[821] <= 16'h7fff;
 filter_in_data_log_force[822] <= 16'h8000;
 filter_in_data_log_force[823] <= 16'h8000;
 filter_in_data_log_force[824] <= 16'h7fff;
 filter_in_data_log_force[825] <= 16'h8000;
 filter_in_data_log_force[826] <= 16'h8000;
 filter_in_data_log_force[827] <= 16'h7fff;
 filter_in_data_log_force[828] <= 16'h7fff;
 filter_in_data_log_force[829] <= 16'h8000;
 filter_in_data_log_force[830] <= 16'h7fff;
 filter_in_data_log_force[831] <= 16'h7fff;
 filter_in_data_log_force[832] <= 16'h8000;
 filter_in_data_log_force[833] <= 16'h7fff;
 filter_in_data_log_force[834] <= 16'h7fff;
 filter_in_data_log_force[835] <= 16'h8000;
 filter_in_data_log_force[836] <= 16'h8000;
 filter_in_data_log_force[837] <= 16'h7fff;
 filter_in_data_log_force[838] <= 16'h8000;
 filter_in_data_log_force[839] <= 16'h8000;
 filter_in_data_log_force[840] <= 16'h7fff;
 filter_in_data_log_force[841] <= 16'h7fff;
 filter_in_data_log_force[842] <= 16'h7fff;
 filter_in_data_log_force[843] <= 16'h7fff;
 filter_in_data_log_force[844] <= 16'h7fff;
 filter_in_data_log_force[845] <= 16'h8000;
 filter_in_data_log_force[846] <= 16'h8000;
 filter_in_data_log_force[847] <= 16'h8000;
 filter_in_data_log_force[848] <= 16'h8000;
 filter_in_data_log_force[849] <= 16'h8000;
 filter_in_data_log_force[850] <= 16'h7fff;
 filter_in_data_log_force[851] <= 16'h8000;
 filter_in_data_log_force[852] <= 16'h8000;
 filter_in_data_log_force[853] <= 16'h7fff;
 filter_in_data_log_force[854] <= 16'h0cee;
 filter_in_data_log_force[855] <= 16'h8000;
 filter_in_data_log_force[856] <= 16'h7fff;
 filter_in_data_log_force[857] <= 16'h7fff;
 filter_in_data_log_force[858] <= 16'h8000;
 filter_in_data_log_force[859] <= 16'h8000;
 filter_in_data_log_force[860] <= 16'h7fff;
 filter_in_data_log_force[861] <= 16'h8000;
 filter_in_data_log_force[862] <= 16'h8000;
 filter_in_data_log_force[863] <= 16'h7fff;
 filter_in_data_log_force[864] <= 16'h7fff;
 filter_in_data_log_force[865] <= 16'h8000;
 filter_in_data_log_force[866] <= 16'h7fff;
 filter_in_data_log_force[867] <= 16'h7fff;
 filter_in_data_log_force[868] <= 16'h7fff;
 filter_in_data_log_force[869] <= 16'h7fff;
 filter_in_data_log_force[870] <= 16'h7fff;
 filter_in_data_log_force[871] <= 16'h7fff;
 filter_in_data_log_force[872] <= 16'h7fff;
 filter_in_data_log_force[873] <= 16'h7fff;
 filter_in_data_log_force[874] <= 16'h7fff;
 filter_in_data_log_force[875] <= 16'h8000;
 filter_in_data_log_force[876] <= 16'h7fff;
 filter_in_data_log_force[877] <= 16'h7fff;
 filter_in_data_log_force[878] <= 16'h8000;
 filter_in_data_log_force[879] <= 16'h7fff;
 filter_in_data_log_force[880] <= 16'h7fff;
 filter_in_data_log_force[881] <= 16'h8000;
 filter_in_data_log_force[882] <= 16'h0000;
 filter_in_data_log_force[883] <= 16'h7fff;
 filter_in_data_log_force[884] <= 16'h8000;
 filter_in_data_log_force[885] <= 16'h8000;
 filter_in_data_log_force[886] <= 16'h7fff;
 filter_in_data_log_force[887] <= 16'h8000;
 filter_in_data_log_force[888] <= 16'h8000;
 filter_in_data_log_force[889] <= 16'h7fff;
 filter_in_data_log_force[890] <= 16'h7fff;
 filter_in_data_log_force[891] <= 16'h8000;
 filter_in_data_log_force[892] <= 16'h7fff;
 filter_in_data_log_force[893] <= 16'h7fff;
 filter_in_data_log_force[894] <= 16'h8000;
 filter_in_data_log_force[895] <= 16'h8000;
 filter_in_data_log_force[896] <= 16'h7fff;
 filter_in_data_log_force[897] <= 16'h8000;
 filter_in_data_log_force[898] <= 16'h8000;
 filter_in_data_log_force[899] <= 16'h7fff;
 filter_in_data_log_force[900] <= 16'h8000;
 filter_in_data_log_force[901] <= 16'h8000;
 filter_in_data_log_force[902] <= 16'h7fff;
 filter_in_data_log_force[903] <= 16'h7fff;
 filter_in_data_log_force[904] <= 16'h8000;
 filter_in_data_log_force[905] <= 16'h8000;
 filter_in_data_log_force[906] <= 16'h7fff;
 filter_in_data_log_force[907] <= 16'h8000;
 filter_in_data_log_force[908] <= 16'h8000;
 filter_in_data_log_force[909] <= 16'h7fff;
 filter_in_data_log_force[910] <= 16'h8000;
 filter_in_data_log_force[911] <= 16'h8000;
 filter_in_data_log_force[912] <= 16'h7fff;
 filter_in_data_log_force[913] <= 16'h8000;
 filter_in_data_log_force[914] <= 16'h8000;
 filter_in_data_log_force[915] <= 16'h7fff;
 filter_in_data_log_force[916] <= 16'h7fff;
 filter_in_data_log_force[917] <= 16'h8000;
 filter_in_data_log_force[918] <= 16'h8000;
 filter_in_data_log_force[919] <= 16'h7fff;
 filter_in_data_log_force[920] <= 16'h8000;
 filter_in_data_log_force[921] <= 16'h8000;
 filter_in_data_log_force[922] <= 16'h7fff;
 filter_in_data_log_force[923] <= 16'h7fff;
 filter_in_data_log_force[924] <= 16'h8000;
 filter_in_data_log_force[925] <= 16'h7fff;
 filter_in_data_log_force[926] <= 16'h7fff;
 filter_in_data_log_force[927] <= 16'h8000;
 filter_in_data_log_force[928] <= 16'h7fff;
 filter_in_data_log_force[929] <= 16'h26af;
 filter_in_data_log_force[930] <= 16'h8000;
 filter_in_data_log_force[931] <= 16'h8000;
 filter_in_data_log_force[932] <= 16'h7fff;
 filter_in_data_log_force[933] <= 16'h8000;
 filter_in_data_log_force[934] <= 16'h8000;
 filter_in_data_log_force[935] <= 16'h7fff;
 filter_in_data_log_force[936] <= 16'h7fff;
 filter_in_data_log_force[937] <= 16'h7fff;
 filter_in_data_log_force[938] <= 16'h7fff;
 filter_in_data_log_force[939] <= 16'h8000;
 filter_in_data_log_force[940] <= 16'h8000;
 filter_in_data_log_force[941] <= 16'h8000;
 filter_in_data_log_force[942] <= 16'h7fff;
 filter_in_data_log_force[943] <= 16'h8000;
 filter_in_data_log_force[944] <= 16'h8000;
 filter_in_data_log_force[945] <= 16'h7fff;
 filter_in_data_log_force[946] <= 16'h8000;
 filter_in_data_log_force[947] <= 16'h8000;
 filter_in_data_log_force[948] <= 16'h7fff;
 filter_in_data_log_force[949] <= 16'h8000;
 filter_in_data_log_force[950] <= 16'h8000;
 filter_in_data_log_force[951] <= 16'h7fff;
 filter_in_data_log_force[952] <= 16'h7fff;
 filter_in_data_log_force[953] <= 16'h8000;
 filter_in_data_log_force[954] <= 16'h7fff;
 filter_in_data_log_force[955] <= 16'h7fff;
 filter_in_data_log_force[956] <= 16'h8000;
 filter_in_data_log_force[957] <= 16'h8000;
 filter_in_data_log_force[958] <= 16'h7fff;
 filter_in_data_log_force[959] <= 16'h7fff;
 filter_in_data_log_force[960] <= 16'h5970;
 filter_in_data_log_force[961] <= 16'h7fff;
 filter_in_data_log_force[962] <= 16'h7fff;
 filter_in_data_log_force[963] <= 16'h8000;
 filter_in_data_log_force[964] <= 16'h7fff;
 filter_in_data_log_force[965] <= 16'h7fff;
 filter_in_data_log_force[966] <= 16'h8000;
 filter_in_data_log_force[967] <= 16'h7fff;
 filter_in_data_log_force[968] <= 16'h7fff;
 filter_in_data_log_force[969] <= 16'h8000;
 filter_in_data_log_force[970] <= 16'h8000;
 filter_in_data_log_force[971] <= 16'h7fff;
 filter_in_data_log_force[972] <= 16'h0000;
 filter_in_data_log_force[973] <= 16'h8000;
 filter_in_data_log_force[974] <= 16'h7fff;
 filter_in_data_log_force[975] <= 16'h7fff;
 filter_in_data_log_force[976] <= 16'h8000;
 filter_in_data_log_force[977] <= 16'h7fff;
 filter_in_data_log_force[978] <= 16'h7fff;
 filter_in_data_log_force[979] <= 16'h8000;
 filter_in_data_log_force[980] <= 16'h8000;
 filter_in_data_log_force[981] <= 16'h7fff;
 filter_in_data_log_force[982] <= 16'h8000;
 filter_in_data_log_force[983] <= 16'h8000;
 filter_in_data_log_force[984] <= 16'h7fff;
 filter_in_data_log_force[985] <= 16'h7fff;
 filter_in_data_log_force[986] <= 16'h8000;
 filter_in_data_log_force[987] <= 16'h7fff;
 filter_in_data_log_force[988] <= 16'h7fff;
 filter_in_data_log_force[989] <= 16'h8000;
 filter_in_data_log_force[990] <= 16'h8000;
 filter_in_data_log_force[991] <= 16'h7fff;
 filter_in_data_log_force[992] <= 16'h8000;
 filter_in_data_log_force[993] <= 16'h8000;
 filter_in_data_log_force[994] <= 16'h7fff;
 filter_in_data_log_force[995] <= 16'h8000;
 filter_in_data_log_force[996] <= 16'h8000;
 filter_in_data_log_force[997] <= 16'h7fff;
 filter_in_data_log_force[998] <= 16'h7fff;
 filter_in_data_log_force[999] <= 16'h8000;

 // Output data for filter_out
 filter_out_expected[  0] <= 12'hffb;
 filter_out_expected[  1] <= 12'hff6;
 filter_out_expected[  2] <= 12'hff4;
 filter_out_expected[  3] <= 12'hffe;
 filter_out_expected[  4] <= 12'h035;
 filter_out_expected[  5] <= 12'h045;
 filter_out_expected[  6] <= 12'hfd8;
 filter_out_expected[  7] <= 12'hfbb;
 filter_out_expected[  8] <= 12'h035;
 filter_out_expected[  9] <= 12'h014;
 filter_out_expected[ 10] <= 12'hfae;
 filter_out_expected[ 11] <= 12'h016;
 filter_out_expected[ 12] <= 12'h019;
 filter_out_expected[ 13] <= 12'hf9b;
 filter_out_expected[ 14] <= 12'h012;
 filter_out_expected[ 15] <= 12'h026;
 filter_out_expected[ 16] <= 12'hf9b;
 filter_out_expected[ 17] <= 12'h03e;
 filter_out_expected[ 18] <= 12'h057;
 filter_out_expected[ 19] <= 12'hfaa;
 filter_out_expected[ 20] <= 12'h021;
 filter_out_expected[ 21] <= 12'h062;
 filter_out_expected[ 22] <= 12'h05f;
 filter_out_expected[ 23] <= 12'h07c;
 filter_out_expected[ 24] <= 12'h0ea;
 filter_out_expected[ 25] <= 12'h09e;
 filter_out_expected[ 26] <= 12'h9b8;
 filter_out_expected[ 27] <= 12'h8d9;
 filter_out_expected[ 28] <= 12'h9be;
 filter_out_expected[ 29] <= 12'hac7;
 filter_out_expected[ 30] <= 12'h75e;
 filter_out_expected[ 31] <= 12'hccf;
 filter_out_expected[ 32] <= 12'h7e8;
 filter_out_expected[ 33] <= 12'ha0c;
 filter_out_expected[ 34] <= 12'hbaa;
 filter_out_expected[ 35] <= 12'h7ee;
 filter_out_expected[ 36] <= 12'hb8d;
 filter_out_expected[ 37] <= 12'ha33;
 filter_out_expected[ 38] <= 12'h850;
 filter_out_expected[ 39] <= 12'hd92;
 filter_out_expected[ 40] <= 12'h75b;
 filter_out_expected[ 41] <= 12'hb46;
 filter_out_expected[ 42] <= 12'ha68;
 filter_out_expected[ 43] <= 12'h6cd;
 filter_out_expected[ 44] <= 12'hcb1;
 filter_out_expected[ 45] <= 12'h6d8;
 filter_out_expected[ 46] <= 12'ha0c;
 filter_out_expected[ 47] <= 12'h9d8;
 filter_out_expected[ 48] <= 12'h6d7;
 filter_out_expected[ 49] <= 12'hb2b;
 filter_out_expected[ 50] <= 12'h5ac;
 filter_out_expected[ 51] <= 12'ha47;
 filter_out_expected[ 52] <= 12'h705;
 filter_out_expected[ 53] <= 12'h946;
 filter_out_expected[ 54] <= 12'h7f4;
 filter_out_expected[ 55] <= 12'h93b;
 filter_out_expected[ 56] <= 12'h690;
 filter_out_expected[ 57] <= 12'hbd8;
 filter_out_expected[ 58] <= 12'h574;
 filter_out_expected[ 59] <= 12'hcb3;
 filter_out_expected[ 60] <= 12'h7be;
 filter_out_expected[ 61] <= 12'h9cc;
 filter_out_expected[ 62] <= 12'hcf5;
 filter_out_expected[ 63] <= 12'h659;
 filter_out_expected[ 64] <= 12'he60;
 filter_out_expected[ 65] <= 12'h8bf;
 filter_out_expected[ 66] <= 12'hc4e;
 filter_out_expected[ 67] <= 12'ha9c;
 filter_out_expected[ 68] <= 12'hce4;
 filter_out_expected[ 69] <= 12'h872;
 filter_out_expected[ 70] <= 12'hed2;
 filter_out_expected[ 71] <= 12'h78b;
 filter_out_expected[ 72] <= 12'hccd;
 filter_out_expected[ 73] <= 12'hb56;
 filter_out_expected[ 74] <= 12'h7bb;
 filter_out_expected[ 75] <= 12'he73;
 filter_out_expected[ 76] <= 12'h76f;
 filter_out_expected[ 77] <= 12'hacf;
 filter_out_expected[ 78] <= 12'hbb0;
 filter_out_expected[ 79] <= 12'h6de;
 filter_out_expected[ 80] <= 12'hbc5;
 filter_out_expected[ 81] <= 12'h71c;
 filter_out_expected[ 82] <= 12'h8c2;
 filter_out_expected[ 83] <= 12'h725;
 filter_out_expected[ 84] <= 12'h8e7;
 filter_out_expected[ 85] <= 12'h325;
 filter_out_expected[ 86] <= 12'h8ad;
 filter_out_expected[ 87] <= 12'h3b2;
 filter_out_expected[ 88] <= 12'h381;
 filter_out_expected[ 89] <= 12'h7b3;
 filter_out_expected[ 90] <= 12'he69;
 filter_out_expected[ 91] <= 12'h71b;
 filter_out_expected[ 92] <= 12'h098;
 filter_out_expected[ 93] <= 12'h074;
 filter_out_expected[ 94] <= 12'h71d;
 filter_out_expected[ 95] <= 12'hda6;
 filter_out_expected[ 96] <= 12'h672;
 filter_out_expected[ 97] <= 12'h358;
 filter_out_expected[ 98] <= 12'h27e;
 filter_out_expected[ 99] <= 12'h7bb;
 filter_out_expected[100] <= 12'h3d2;
 filter_out_expected[101] <= 12'h663;
 filter_out_expected[102] <= 12'h8d1;
 filter_out_expected[103] <= 12'h463;
 filter_out_expected[104] <= 12'ha4d;
 filter_out_expected[105] <= 12'h5ce;
 filter_out_expected[106] <= 12'h919;
 filter_out_expected[107] <= 12'h72f;
 filter_out_expected[108] <= 12'h968;
 filter_out_expected[109] <= 12'h6a8;
 filter_out_expected[110] <= 12'ha59;
 filter_out_expected[111] <= 12'h698;
 filter_out_expected[112] <= 12'ha2b;
 filter_out_expected[113] <= 12'h752;
 filter_out_expected[114] <= 12'h9e9;
 filter_out_expected[115] <= 12'h6ae;
 filter_out_expected[116] <= 12'haf9;
 filter_out_expected[117] <= 12'h6b9;
 filter_out_expected[118] <= 12'h992;
 filter_out_expected[119] <= 12'h940;
 filter_out_expected[120] <= 12'h6d3;
 filter_out_expected[121] <= 12'hb0f;
 filter_out_expected[122] <= 12'h626;
 filter_out_expected[123] <= 12'ha64;
 filter_out_expected[124] <= 12'h753;
 filter_out_expected[125] <= 12'h96d;
 filter_out_expected[126] <= 12'h783;
 filter_out_expected[127] <= 12'habf;
 filter_out_expected[128] <= 12'h6eb;
 filter_out_expected[129] <= 12'hb39;
 filter_out_expected[130] <= 12'h6b3;
 filter_out_expected[131] <= 12'h956;
 filter_out_expected[132] <= 12'h894;
 filter_out_expected[133] <= 12'h638;
 filter_out_expected[134] <= 12'hb38;
 filter_out_expected[135] <= 12'h5b0;
 filter_out_expected[136] <= 12'h9d4;
 filter_out_expected[137] <= 12'h75f;
 filter_out_expected[138] <= 12'h902;
 filter_out_expected[139] <= 12'h79f;
 filter_out_expected[140] <= 12'hab7;
 filter_out_expected[141] <= 12'h637;
 filter_out_expected[142] <= 12'hc4a;
 filter_out_expected[143] <= 12'h7d2;
 filter_out_expected[144] <= 12'ha99;
 filter_out_expected[145] <= 12'hbe8;
 filter_out_expected[146] <= 12'h7e1;
 filter_out_expected[147] <= 12'he6a;
 filter_out_expected[148] <= 12'h7f8;
 filter_out_expected[149] <= 12'hd00;
 filter_out_expected[150] <= 12'ha06;
 filter_out_expected[151] <= 12'hc1f;
 filter_out_expected[152] <= 12'h8f7;
 filter_out_expected[153] <= 12'hdd2;
 filter_out_expected[154] <= 12'h71d;
 filter_out_expected[155] <= 12'hdad;
 filter_out_expected[156] <= 12'h93c;
 filter_out_expected[157] <= 12'ha2e;
 filter_out_expected[158] <= 12'he5d;
 filter_out_expected[159] <= 12'h59d;
 filter_out_expected[160] <= 12'h1cd;
 filter_out_expected[161] <= 12'h622;
 filter_out_expected[162] <= 12'hf8f;
 filter_out_expected[163] <= 12'ha1b;
 filter_out_expected[164] <= 12'hba2;
 filter_out_expected[165] <= 12'hbf0;
 filter_out_expected[166] <= 12'h998;
 filter_out_expected[167] <= 12'hb6f;
 filter_out_expected[168] <= 12'h6dc;
 filter_out_expected[169] <= 12'haee;
 filter_out_expected[170] <= 12'h435;
 filter_out_expected[171] <= 12'h820;
 filter_out_expected[172] <= 12'h4a3;
 filter_out_expected[173] <= 12'h1d8;
 filter_out_expected[174] <= 12'h5a0;
 filter_out_expected[175] <= 12'hdf6;
 filter_out_expected[176] <= 12'h3f5;
 filter_out_expected[177] <= 12'hf9d;
 filter_out_expected[178] <= 12'h095;
 filter_out_expected[179] <= 12'h265;
 filter_out_expected[180] <= 12'h054;
 filter_out_expected[181] <= 12'h0fb;
 filter_out_expected[182] <= 12'h55f;
 filter_out_expected[183] <= 12'h075;
 filter_out_expected[184] <= 12'h84d;
 filter_out_expected[185] <= 12'h38b;
 filter_out_expected[186] <= 12'h87f;
 filter_out_expected[187] <= 12'h689;
 filter_out_expected[188] <= 12'h9f1;
 filter_out_expected[189] <= 12'h7ea;
 filter_out_expected[190] <= 12'ha96;
 filter_out_expected[191] <= 12'h96f;
 filter_out_expected[192] <= 12'h85a;
 filter_out_expected[193] <= 12'hbd9;
 filter_out_expected[194] <= 12'h673;
 filter_out_expected[195] <= 12'hb58;
 filter_out_expected[196] <= 12'h727;
 filter_out_expected[197] <= 12'h946;
 filter_out_expected[198] <= 12'h7ae;
 filter_out_expected[199] <= 12'h927;
 filter_out_expected[200] <= 12'h5c5;
 filter_out_expected[201] <= 12'hb35;
 filter_out_expected[202] <= 12'h5b2;
 filter_out_expected[203] <= 12'h97f;
 filter_out_expected[204] <= 12'h9e5;
 filter_out_expected[205] <= 12'h6b2;
 filter_out_expected[206] <= 12'hcfc;
 filter_out_expected[207] <= 12'h72b;
 filter_out_expected[208] <= 12'hae0;
 filter_out_expected[209] <= 12'hba9;
 filter_out_expected[210] <= 12'h7ac;
 filter_out_expected[211] <= 12'hdcf;
 filter_out_expected[212] <= 12'h897;
 filter_out_expected[213] <= 12'ha9f;
 filter_out_expected[214] <= 12'hb33;
 filter_out_expected[215] <= 12'h752;
 filter_out_expected[216] <= 12'hb21;
 filter_out_expected[217] <= 12'h8b8;
 filter_out_expected[218] <= 12'h732;
 filter_out_expected[219] <= 12'hbd6;
 filter_out_expected[220] <= 12'h59f;
 filter_out_expected[221] <= 12'haa8;
 filter_out_expected[222] <= 12'h756;
 filter_out_expected[223] <= 12'h914;
 filter_out_expected[224] <= 12'h80d;
 filter_out_expected[225] <= 12'ha0a;
 filter_out_expected[226] <= 12'h639;
 filter_out_expected[227] <= 12'hbb7;
 filter_out_expected[228] <= 12'h648;
 filter_out_expected[229] <= 12'ha31;
 filter_out_expected[230] <= 12'h9bb;
 filter_out_expected[231] <= 12'h5a8;
 filter_out_expected[232] <= 12'hdcc;
 filter_out_expected[233] <= 12'h39c;
 filter_out_expected[234] <= 12'hcec;
 filter_out_expected[235] <= 12'h6bd;
 filter_out_expected[236] <= 12'h8a5;
 filter_out_expected[237] <= 12'hb16;
 filter_out_expected[238] <= 12'h6fc;
 filter_out_expected[239] <= 12'hbe4;
 filter_out_expected[240] <= 12'h8cf;
 filter_out_expected[241] <= 12'hb71;
 filter_out_expected[242] <= 12'ha20;
 filter_out_expected[243] <= 12'he0b;
 filter_out_expected[244] <= 12'h79d;
 filter_out_expected[245] <= 12'h240;
 filter_out_expected[246] <= 12'h6af;
 filter_out_expected[247] <= 12'h0f7;
 filter_out_expected[248] <= 12'ha35;
 filter_out_expected[249] <= 12'hc02;
 filter_out_expected[250] <= 12'hc74;
 filter_out_expected[251] <= 12'h914;
 filter_out_expected[252] <= 12'hb59;
 filter_out_expected[253] <= 12'h6b3;
 filter_out_expected[254] <= 12'ha14;
 filter_out_expected[255] <= 12'h413;
 filter_out_expected[256] <= 12'h7e7;
 filter_out_expected[257] <= 12'h3cf;
 filter_out_expected[258] <= 12'h20a;
 filter_out_expected[259] <= 12'h5fc;
 filter_out_expected[260] <= 12'he49;
 filter_out_expected[261] <= 12'h5a1;
 filter_out_expected[262] <= 12'h035;
 filter_out_expected[263] <= 12'h0db;
 filter_out_expected[264] <= 12'h50d;
 filter_out_expected[265] <= 12'hee5;
 filter_out_expected[266] <= 12'ha8d;
 filter_out_expected[267] <= 12'h3fa;
 filter_out_expected[268] <= 12'h314;
 filter_out_expected[269] <= 12'h89e;
 filter_out_expected[270] <= 12'h413;
 filter_out_expected[271] <= 12'h99f;
 filter_out_expected[272] <= 12'h681;
 filter_out_expected[273] <= 12'ha58;
 filter_out_expected[274] <= 12'h833;
 filter_out_expected[275] <= 12'ha5d;
 filter_out_expected[276] <= 12'h9a0;
 filter_out_expected[277] <= 12'h83b;
 filter_out_expected[278] <= 12'hbd1;
 filter_out_expected[279] <= 12'h69d;
 filter_out_expected[280] <= 12'hb4a;
 filter_out_expected[281] <= 12'h79b;
 filter_out_expected[282] <= 12'h8a5;
 filter_out_expected[283] <= 12'h5c5;
 filter_out_expected[284] <= 12'h8e5;
 filter_out_expected[285] <= 12'h655;
 filter_out_expected[286] <= 12'hb39;
 filter_out_expected[287] <= 12'h647;
 filter_out_expected[288] <= 12'ha03;
 filter_out_expected[289] <= 12'ha2a;
 filter_out_expected[290] <= 12'h71b;
 filter_out_expected[291] <= 12'hd06;
 filter_out_expected[292] <= 12'h778;
 filter_out_expected[293] <= 12'hb24;
 filter_out_expected[294] <= 12'hbbf;
 filter_out_expected[295] <= 12'h83a;
 filter_out_expected[296] <= 12'hd20;
 filter_out_expected[297] <= 12'h787;
 filter_out_expected[298] <= 12'ha34;
 filter_out_expected[299] <= 12'h92e;
 filter_out_expected[300] <= 12'h691;
 filter_out_expected[301] <= 12'hafd;
 filter_out_expected[302] <= 12'h4e5;
 filter_out_expected[303] <= 12'h94f;
 filter_out_expected[304] <= 12'h5ee;
 filter_out_expected[305] <= 12'h7d7;
 filter_out_expected[306] <= 12'h6f0;
 filter_out_expected[307] <= 12'h826;
 filter_out_expected[308] <= 12'h775;
 filter_out_expected[309] <= 12'h2cf;
 filter_out_expected[310] <= 12'h968;
 filter_out_expected[311] <= 12'h7c5;
 filter_out_expected[312] <= 12'hbaf;
 filter_out_expected[313] <= 12'h795;
 filter_out_expected[314] <= 12'hd2e;
 filter_out_expected[315] <= 12'h836;
 filter_out_expected[316] <= 12'hcc7;
 filter_out_expected[317] <= 12'h988;
 filter_out_expected[318] <= 12'hc9a;
 filter_out_expected[319] <= 12'h8e1;
 filter_out_expected[320] <= 12'hdbb;
 filter_out_expected[321] <= 12'h78b;
 filter_out_expected[322] <= 12'hd61;
 filter_out_expected[323] <= 12'h91d;
 filter_out_expected[324] <= 12'ha5f;
 filter_out_expected[325] <= 12'hdc4;
 filter_out_expected[326] <= 12'h591;
 filter_out_expected[327] <= 12'h1f2;
 filter_out_expected[328] <= 12'h58b;
 filter_out_expected[329] <= 12'h036;
 filter_out_expected[330] <= 12'ha99;
 filter_out_expected[331] <= 12'hb80;
 filter_out_expected[332] <= 12'hdcf;
 filter_out_expected[333] <= 12'ha23;
 filter_out_expected[334] <= 12'hbd7;
 filter_out_expected[335] <= 12'hb14;
 filter_out_expected[336] <= 12'h89b;
 filter_out_expected[337] <= 12'ha5b;
 filter_out_expected[338] <= 12'h62d;
 filter_out_expected[339] <= 12'h8aa;
 filter_out_expected[340] <= 12'h2ba;
 filter_out_expected[341] <= 12'h6d9;
 filter_out_expected[342] <= 12'hfdf;
 filter_out_expected[343] <= 12'h47f;
 filter_out_expected[344] <= 12'h067;
 filter_out_expected[345] <= 12'h0fd;
 filter_out_expected[346] <= 12'h25c;
 filter_out_expected[347] <= 12'hfef;
 filter_out_expected[348] <= 12'h02b;
 filter_out_expected[349] <= 12'h4c3;
 filter_out_expected[350] <= 12'he8a;
 filter_out_expected[351] <= 12'h700;
 filter_out_expected[352] <= 12'h28c;
 filter_out_expected[353] <= 12'h47a;
 filter_out_expected[354] <= 12'h8bb;
 filter_out_expected[355] <= 12'h413;
 filter_out_expected[356] <= 12'ha3d;
 filter_out_expected[357] <= 12'h68e;
 filter_out_expected[358] <= 12'h95e;
 filter_out_expected[359] <= 12'h7c7;
 filter_out_expected[360] <= 12'ha22;
 filter_out_expected[361] <= 12'h6b7;
 filter_out_expected[362] <= 12'ha07;
 filter_out_expected[363] <= 12'h4fe;
 filter_out_expected[364] <= 12'h8da;
 filter_out_expected[365] <= 12'h7fe;
 filter_out_expected[366] <= 12'h995;
 filter_out_expected[367] <= 12'h5fb;
 filter_out_expected[368] <= 12'hc12;
 filter_out_expected[369] <= 12'h6a1;
 filter_out_expected[370] <= 12'h9e4;
 filter_out_expected[371] <= 12'hbca;
 filter_out_expected[372] <= 12'h7a6;
 filter_out_expected[373] <= 12'hd92;
 filter_out_expected[374] <= 12'hb14;
 filter_out_expected[375] <= 12'h8c2;
 filter_out_expected[376] <= 12'h1ad;
 filter_out_expected[377] <= 12'h538;
 filter_out_expected[378] <= 12'h1de;
 filter_out_expected[379] <= 12'h8e7;
 filter_out_expected[380] <= 12'hb35;
 filter_out_expected[381] <= 12'hd1c;
 filter_out_expected[382] <= 12'h736;
 filter_out_expected[383] <= 12'hc0c;
 filter_out_expected[384] <= 12'h9cf;
 filter_out_expected[385] <= 12'h69e;
 filter_out_expected[386] <= 12'hc22;
 filter_out_expected[387] <= 12'h599;
 filter_out_expected[388] <= 12'h9fb;
 filter_out_expected[389] <= 12'h7c6;
 filter_out_expected[390] <= 12'h897;
 filter_out_expected[391] <= 12'h774;
 filter_out_expected[392] <= 12'ha81;
 filter_out_expected[393] <= 12'h533;
 filter_out_expected[394] <= 12'hb52;
 filter_out_expected[395] <= 12'h69e;
 filter_out_expected[396] <= 12'h850;
 filter_out_expected[397] <= 12'h9da;
 filter_out_expected[398] <= 12'h5d6;
 filter_out_expected[399] <= 12'ha2a;
 filter_out_expected[400] <= 12'h6ff;
 filter_out_expected[401] <= 12'h6f2;
 filter_out_expected[402] <= 12'h971;
 filter_out_expected[403] <= 12'h6c6;
 filter_out_expected[404] <= 12'h788;
 filter_out_expected[405] <= 12'hbc2;
 filter_out_expected[406] <= 12'h3c2;
 filter_out_expected[407] <= 12'hf0f;
 filter_out_expected[408] <= 12'h541;
 filter_out_expected[409] <= 12'hc83;
 filter_out_expected[410] <= 12'hc49;
 filter_out_expected[411] <= 12'h6ff;
 filter_out_expected[412] <= 12'h244;
 filter_out_expected[413] <= 12'h5e5;
 filter_out_expected[414] <= 12'h090;
 filter_out_expected[415] <= 12'ha24;
 filter_out_expected[416] <= 12'hb7f;
 filter_out_expected[417] <= 12'hc54;
 filter_out_expected[418] <= 12'h906;
 filter_out_expected[419] <= 12'hb09;
 filter_out_expected[420] <= 12'h6c8;
 filter_out_expected[421] <= 12'ha0c;
 filter_out_expected[422] <= 12'h3f3;
 filter_out_expected[423] <= 12'h7f3;
 filter_out_expected[424] <= 12'h3c1;
 filter_out_expected[425] <= 12'h273;
 filter_out_expected[426] <= 12'h66d;
 filter_out_expected[427] <= 12'he7a;
 filter_out_expected[428] <= 12'h652;
 filter_out_expected[429] <= 12'h02e;
 filter_out_expected[430] <= 12'h0b4;
 filter_out_expected[431] <= 12'h66d;
 filter_out_expected[432] <= 12'he39;
 filter_out_expected[433] <= 12'h731;
 filter_out_expected[434] <= 12'h340;
 filter_out_expected[435] <= 12'h48f;
 filter_out_expected[436] <= 12'h8e1;
 filter_out_expected[437] <= 12'h45d;
 filter_out_expected[438] <= 12'ha5d;
 filter_out_expected[439] <= 12'h688;
 filter_out_expected[440] <= 12'ha86;
 filter_out_expected[441] <= 12'h879;
 filter_out_expected[442] <= 12'ha1c;
 filter_out_expected[443] <= 12'h996;
 filter_out_expected[444] <= 12'h82b;
 filter_out_expected[445] <= 12'hb4b;
 filter_out_expected[446] <= 12'h671;
 filter_out_expected[447] <= 12'hafd;
 filter_out_expected[448] <= 12'h6d9;
 filter_out_expected[449] <= 12'h956;
 filter_out_expected[450] <= 12'h777;
 filter_out_expected[451] <= 12'h92b;
 filter_out_expected[452] <= 12'h5f0;
 filter_out_expected[453] <= 12'hb1e;
 filter_out_expected[454] <= 12'h5e4;
 filter_out_expected[455] <= 12'h9d3;
 filter_out_expected[456] <= 12'h9e4;
 filter_out_expected[457] <= 12'h69c;
 filter_out_expected[458] <= 12'hcf2;
 filter_out_expected[459] <= 12'h722;
 filter_out_expected[460] <= 12'hae0;
 filter_out_expected[461] <= 12'hba1;
 filter_out_expected[462] <= 12'h799;
 filter_out_expected[463] <= 12'hdaf;
 filter_out_expected[464] <= 12'h881;
 filter_out_expected[465] <= 12'hafc;
 filter_out_expected[466] <= 12'hbc4;
 filter_out_expected[467] <= 12'h784;
 filter_out_expected[468] <= 12'hb35;
 filter_out_expected[469] <= 12'h893;
 filter_out_expected[470] <= 12'h6cd;
 filter_out_expected[471] <= 12'hbc6;
 filter_out_expected[472] <= 12'h537;
 filter_out_expected[473] <= 12'h9fb;
 filter_out_expected[474] <= 12'h730;
 filter_out_expected[475] <= 12'h873;
 filter_out_expected[476] <= 12'h79d;
 filter_out_expected[477] <= 12'ha5d;
 filter_out_expected[478] <= 12'h5e9;
 filter_out_expected[479] <= 12'hc5a;
 filter_out_expected[480] <= 12'h79b;
 filter_out_expected[481] <= 12'ha9d;
 filter_out_expected[482] <= 12'hc13;
 filter_out_expected[483] <= 12'h7ca;
 filter_out_expected[484] <= 12'he9d;
 filter_out_expected[485] <= 12'h84c;
 filter_out_expected[486] <= 12'hd00;
 filter_out_expected[487] <= 12'h9f0;
 filter_out_expected[488] <= 12'hc15;
 filter_out_expected[489] <= 12'h8ee;
 filter_out_expected[490] <= 12'hdd2;
 filter_out_expected[491] <= 12'h71d;
 filter_out_expected[492] <= 12'hdad;
 filter_out_expected[493] <= 12'h93c;
 filter_out_expected[494] <= 12'ha2e;
 filter_out_expected[495] <= 12'he5d;
 filter_out_expected[496] <= 12'h59d;
 filter_out_expected[497] <= 12'h1cd;
 filter_out_expected[498] <= 12'h622;
 filter_out_expected[499] <= 12'hf8f;
 filter_out_expected[500] <= 12'ha1b;
 filter_out_expected[501] <= 12'hba2;
 filter_out_expected[502] <= 12'hbf0;
 filter_out_expected[503] <= 12'h998;
 filter_out_expected[504] <= 12'hb78;
 filter_out_expected[505] <= 12'h6e7;
 filter_out_expected[506] <= 12'hb04;
 filter_out_expected[507] <= 12'h435;
 filter_out_expected[508] <= 12'h7cc;
 filter_out_expected[509] <= 12'h470;
 filter_out_expected[510] <= 12'h1ef;
 filter_out_expected[511] <= 12'h575;
 filter_out_expected[512] <= 12'hdf1;
 filter_out_expected[513] <= 12'h42b;
 filter_out_expected[514] <= 12'hf8c;
 filter_out_expected[515] <= 12'h0e3;
 filter_out_expected[516] <= 12'h2c0;
 filter_out_expected[517] <= 12'h060;
 filter_out_expected[518] <= 12'h194;
 filter_out_expected[519] <= 12'h5a5;
 filter_out_expected[520] <= 12'h04e;
 filter_out_expected[521] <= 12'h872;
 filter_out_expected[522] <= 12'h2ca;
 filter_out_expected[523] <= 12'h801;
 filter_out_expected[524] <= 12'h65e;
 filter_out_expected[525] <= 12'h80e;
 filter_out_expected[526] <= 12'h74f;
 filter_out_expected[527] <= 12'h9f1;
 filter_out_expected[528] <= 12'h5a2;
 filter_out_expected[529] <= 12'hadd;
 filter_out_expected[530] <= 12'h5b8;
 filter_out_expected[531] <= 12'h934;
 filter_out_expected[532] <= 12'h783;
 filter_out_expected[533] <= 12'h66c;
 filter_out_expected[534] <= 12'h89b;
 filter_out_expected[535] <= 12'h505;
 filter_out_expected[536] <= 12'h8a0;
 filter_out_expected[537] <= 12'h4f0;
 filter_out_expected[538] <= 12'h8c3;
 filter_out_expected[539] <= 12'h5e5;
 filter_out_expected[540] <= 12'h8e6;
 filter_out_expected[541] <= 12'h630;
 filter_out_expected[542] <= 12'h9ee;
 filter_out_expected[543] <= 12'h6e2;
 filter_out_expected[544] <= 12'ha11;
 filter_out_expected[545] <= 12'h772;
 filter_out_expected[546] <= 12'ha9b;
 filter_out_expected[547] <= 12'h6ea;
 filter_out_expected[548] <= 12'hb16;
 filter_out_expected[549] <= 12'h6ed;
 filter_out_expected[550] <= 12'h97f;
 filter_out_expected[551] <= 12'h921;
 filter_out_expected[552] <= 12'h6c9;
 filter_out_expected[553] <= 12'hb06;
 filter_out_expected[554] <= 12'h626;
 filter_out_expected[555] <= 12'ha64;
 filter_out_expected[556] <= 12'h75c;
 filter_out_expected[557] <= 12'h981;
 filter_out_expected[558] <= 12'h7a4;
 filter_out_expected[559] <= 12'had6;
 filter_out_expected[560] <= 12'h68f;
 filter_out_expected[561] <= 12'haa8;
 filter_out_expected[562] <= 12'h681;
 filter_out_expected[563] <= 12'h942;
 filter_out_expected[564] <= 12'h8b9;
 filter_out_expected[565] <= 12'h69e;
 filter_out_expected[566] <= 12'hb47;
 filter_out_expected[567] <= 12'h619;
 filter_out_expected[568] <= 12'ha81;
 filter_out_expected[569] <= 12'h786;
 filter_out_expected[570] <= 12'h9a3;
 filter_out_expected[571] <= 12'h80f;
 filter_out_expected[572] <= 12'ha65;
 filter_out_expected[573] <= 12'h687;
 filter_out_expected[574] <= 12'hba7;
 filter_out_expected[575] <= 12'h67f;
 filter_out_expected[576] <= 12'ha2c;
 filter_out_expected[577] <= 12'h990;
 filter_out_expected[578] <= 12'h5c0;
 filter_out_expected[579] <= 12'hd99;
 filter_out_expected[580] <= 12'h348;
 filter_out_expected[581] <= 12'hcec;
 filter_out_expected[582] <= 12'h6d3;
 filter_out_expected[583] <= 12'h8af;
 filter_out_expected[584] <= 12'hb1f;
 filter_out_expected[585] <= 12'h6fc;
 filter_out_expected[586] <= 12'hbe4;
 filter_out_expected[587] <= 12'h8d5;
 filter_out_expected[588] <= 12'hb78;
 filter_out_expected[589] <= 12'ha2e;
 filter_out_expected[590] <= 12'he0b;
 filter_out_expected[591] <= 12'h767;
 filter_out_expected[592] <= 12'h21f;
 filter_out_expected[593] <= 12'h6be;
 filter_out_expected[594] <= 12'h0e4;
 filter_out_expected[595] <= 12'ha3d;
 filter_out_expected[596] <= 12'hc3c;
 filter_out_expected[597] <= 12'hc69;
 filter_out_expected[598] <= 12'h8f3;
 filter_out_expected[599] <= 12'hb61;
 filter_out_expected[600] <= 12'h6cc;
 filter_out_expected[601] <= 12'ha46;
 filter_out_expected[602] <= 12'h42d;
 filter_out_expected[603] <= 12'h805;
 filter_out_expected[604] <= 12'h410;
 filter_out_expected[605] <= 12'h1fd;
 filter_out_expected[606] <= 12'h5fa;
 filter_out_expected[607] <= 12'he4b;
 filter_out_expected[608] <= 12'h4eb;
 filter_out_expected[609] <= 12'hfd4;
 filter_out_expected[610] <= 12'h057;
 filter_out_expected[611] <= 12'h2d4;
 filter_out_expected[612] <= 12'hfbd;
 filter_out_expected[613] <= 12'h066;
 filter_out_expected[614] <= 12'h560;
 filter_out_expected[615] <= 12'he96;
 filter_out_expected[616] <= 12'h77b;
 filter_out_expected[617] <= 12'h2f7;
 filter_out_expected[618] <= 12'h464;
 filter_out_expected[619] <= 12'h8b1;
 filter_out_expected[620] <= 12'h3c5;
 filter_out_expected[621] <= 12'ha12;
 filter_out_expected[622] <= 12'h67b;
 filter_out_expected[623] <= 12'h8db;
 filter_out_expected[624] <= 12'h789;
 filter_out_expected[625] <= 12'h9fb;
 filter_out_expected[626] <= 12'h674;
 filter_out_expected[627] <= 12'hac3;
 filter_out_expected[628] <= 12'h698;
 filter_out_expected[629] <= 12'h9c0;
 filter_out_expected[630] <= 12'h77e;
 filter_out_expected[631] <= 12'h94b;
 filter_out_expected[632] <= 12'h63d;
 filter_out_expected[633] <= 12'hb37;
 filter_out_expected[634] <= 12'h660;
 filter_out_expected[635] <= 12'ha00;
 filter_out_expected[636] <= 12'h9bd;
 filter_out_expected[637] <= 12'h713;
 filter_out_expected[638] <= 12'hd05;
 filter_out_expected[639] <= 12'h6d4;
 filter_out_expected[640] <= 12'hb27;
 filter_out_expected[641] <= 12'hb33;
 filter_out_expected[642] <= 12'h6b7;
 filter_out_expected[643] <= 12'hd90;
 filter_out_expected[644] <= 12'h7cc;
 filter_out_expected[645] <= 12'ha1c;
 filter_out_expected[646] <= 12'hbca;
 filter_out_expected[647] <= 12'h720;
 filter_out_expected[648] <= 12'hb8e;
 filter_out_expected[649] <= 12'ha13;
 filter_out_expected[650] <= 12'h777;
 filter_out_expected[651] <= 12'hd70;
 filter_out_expected[652] <= 12'h721;
 filter_out_expected[653] <= 12'hb37;
 filter_out_expected[654] <= 12'hba7;
 filter_out_expected[655] <= 12'h7ca;
 filter_out_expected[656] <= 12'hd27;
 filter_out_expected[657] <= 12'h7d3;
 filter_out_expected[658] <= 12'ha56;
 filter_out_expected[659] <= 12'h92e;
 filter_out_expected[660] <= 12'h65a;
 filter_out_expected[661] <= 12'ha43;
 filter_out_expected[662] <= 12'h46e;
 filter_out_expected[663] <= 12'h938;
 filter_out_expected[664] <= 12'h54c;
 filter_out_expected[665] <= 12'h7e1;
 filter_out_expected[666] <= 12'h6ca;
 filter_out_expected[667] <= 12'h687;
 filter_out_expected[668] <= 12'h8a6;
 filter_out_expected[669] <= 12'h670;
 filter_out_expected[670] <= 12'ha4c;
 filter_out_expected[671] <= 12'h75d;
 filter_out_expected[672] <= 12'hbbe;
 filter_out_expected[673] <= 12'h79d;
 filter_out_expected[674] <= 12'hdc6;
 filter_out_expected[675] <= 12'h7b5;
 filter_out_expected[676] <= 12'hcbb;
 filter_out_expected[677] <= 12'hb1a;
 filter_out_expected[678] <= 12'h871;
 filter_out_expected[679] <= 12'he25;
 filter_out_expected[680] <= 12'h6dd;
 filter_out_expected[681] <= 12'hbc3;
 filter_out_expected[682] <= 12'hb17;
 filter_out_expected[683] <= 12'h6d0;
 filter_out_expected[684] <= 12'he69;
 filter_out_expected[685] <= 12'h712;
 filter_out_expected[686] <= 12'hb04;
 filter_out_expected[687] <= 12'hd70;
 filter_out_expected[688] <= 12'h750;
 filter_out_expected[689] <= 12'h017;
 filter_out_expected[690] <= 12'h9ac;
 filter_out_expected[691] <= 12'hc9c;
 filter_out_expected[692] <= 12'hd90;
 filter_out_expected[693] <= 12'ha3e;
 filter_out_expected[694] <= 12'hd01;
 filter_out_expected[695] <= 12'hac5;
 filter_out_expected[696] <= 12'h977;
 filter_out_expected[697] <= 12'hb6f;
 filter_out_expected[698] <= 12'h608;
 filter_out_expected[699] <= 12'ha99;
 filter_out_expected[700] <= 12'h396;
 filter_out_expected[701] <= 12'h737;
 filter_out_expected[702] <= 12'h3ee;
 filter_out_expected[703] <= 12'h1f2;
 filter_out_expected[704] <= 12'h5ff;
 filter_out_expected[705] <= 12'hea2;
 filter_out_expected[706] <= 12'h67f;
 filter_out_expected[707] <= 12'h0d4;
 filter_out_expected[708] <= 12'h170;
 filter_out_expected[709] <= 12'h6b9;
 filter_out_expected[710] <= 12'he7d;
 filter_out_expected[711] <= 12'h7ab;
 filter_out_expected[712] <= 12'h338;
 filter_out_expected[713] <= 12'h405;
 filter_out_expected[714] <= 12'h8b7;
 filter_out_expected[715] <= 12'h39a;
 filter_out_expected[716] <= 12'h95a;
 filter_out_expected[717] <= 12'h62e;
 filter_out_expected[718] <= 12'h8ca;
 filter_out_expected[719] <= 12'h764;
 filter_out_expected[720] <= 12'ha06;
 filter_out_expected[721] <= 12'h65e;
 filter_out_expected[722] <= 12'haad;
 filter_out_expected[723] <= 12'h708;
 filter_out_expected[724] <= 12'ha03;
 filter_out_expected[725] <= 12'h7b3;
 filter_out_expected[726] <= 12'ha2e;
 filter_out_expected[727] <= 12'h66c;
 filter_out_expected[728] <= 12'hafa;
 filter_out_expected[729] <= 12'h6d0;
 filter_out_expected[730] <= 12'h968;
 filter_out_expected[731] <= 12'h929;
 filter_out_expected[732] <= 12'h714;
 filter_out_expected[733] <= 12'hb26;
 filter_out_expected[734] <= 12'h603;
 filter_out_expected[735] <= 12'ha93;
 filter_out_expected[736] <= 12'h719;
 filter_out_expected[737] <= 12'h8df;
 filter_out_expected[738] <= 12'h764;
 filter_out_expected[739] <= 12'h9f4;
 filter_out_expected[740] <= 12'h601;
 filter_out_expected[741] <= 12'hb36;
 filter_out_expected[742] <= 12'h64f;
 filter_out_expected[743] <= 12'h9af;
 filter_out_expected[744] <= 12'ha13;
 filter_out_expected[745] <= 12'h6ec;
 filter_out_expected[746] <= 12'hceb;
 filter_out_expected[747] <= 12'h7b1;
 filter_out_expected[748] <= 12'hb19;
 filter_out_expected[749] <= 12'hb8d;
 filter_out_expected[750] <= 12'h83c;
 filter_out_expected[751] <= 12'hd41;
 filter_out_expected[752] <= 12'h7a6;
 filter_out_expected[753] <= 12'ha62;
 filter_out_expected[754] <= 12'h955;
 filter_out_expected[755] <= 12'h65f;
 filter_out_expected[756] <= 12'hae7;
 filter_out_expected[757] <= 12'h51e;
 filter_out_expected[758] <= 12'h933;
 filter_out_expected[759] <= 12'h5d7;
 filter_out_expected[760] <= 12'h7fe;
 filter_out_expected[761] <= 12'h686;
 filter_out_expected[762] <= 12'h737;
 filter_out_expected[763] <= 12'h7cc;
 filter_out_expected[764] <= 12'h5b0;
 filter_out_expected[765] <= 12'ha89;
 filter_out_expected[766] <= 12'h4aa;
 filter_out_expected[767] <= 12'habb;
 filter_out_expected[768] <= 12'h723;
 filter_out_expected[769] <= 12'h82f;
 filter_out_expected[770] <= 12'ha25;
 filter_out_expected[771] <= 12'h66b;
 filter_out_expected[772] <= 12'ha2f;
 filter_out_expected[773] <= 12'h7fe;
 filter_out_expected[774] <= 12'h77a;
 filter_out_expected[775] <= 12'h943;
 filter_out_expected[776] <= 12'h777;
 filter_out_expected[777] <= 12'h6f6;
 filter_out_expected[778] <= 12'hb03;
 filter_out_expected[779] <= 12'h3da;
 filter_out_expected[780] <= 12'hcfe;
 filter_out_expected[781] <= 12'h41c;
 filter_out_expected[782] <= 12'hbef;
 filter_out_expected[783] <= 12'h845;
 filter_out_expected[784] <= 12'h931;
 filter_out_expected[785] <= 12'hc21;
 filter_out_expected[786] <= 12'h80e;
 filter_out_expected[787] <= 12'hc75;
 filter_out_expected[788] <= 12'h990;
 filter_out_expected[789] <= 12'haae;
 filter_out_expected[790] <= 12'ha76;
 filter_out_expected[791] <= 12'h907;
 filter_out_expected[792] <= 12'ha75;
 filter_out_expected[793] <= 12'h639;
 filter_out_expected[794] <= 12'ha85;
 filter_out_expected[795] <= 12'h3cc;
 filter_out_expected[796] <= 12'h822;
 filter_out_expected[797] <= 12'h44e;
 filter_out_expected[798] <= 12'h274;
 filter_out_expected[799] <= 12'h6c4;
 filter_out_expected[800] <= 12'hec8;
 filter_out_expected[801] <= 12'h64f;
 filter_out_expected[802] <= 12'h06c;
 filter_out_expected[803] <= 12'h0ac;
 filter_out_expected[804] <= 12'h648;
 filter_out_expected[805] <= 12'he51;
 filter_out_expected[806] <= 12'h6f6;
 filter_out_expected[807] <= 12'h2ee;
 filter_out_expected[808] <= 12'h483;
 filter_out_expected[809] <= 12'h8e8;
 filter_out_expected[810] <= 12'h467;
 filter_out_expected[811] <= 12'ha4f;
 filter_out_expected[812] <= 12'h680;
 filter_out_expected[813] <= 12'ha8c;
 filter_out_expected[814] <= 12'h865;
 filter_out_expected[815] <= 12'ha32;
 filter_out_expected[816] <= 12'h9ad;
 filter_out_expected[817] <= 12'h82b;
 filter_out_expected[818] <= 12'hb9f;
 filter_out_expected[819] <= 12'h69c;
 filter_out_expected[820] <= 12'hb2b;
 filter_out_expected[821] <= 12'h780;
 filter_out_expected[822] <= 12'h8ab;
 filter_out_expected[823] <= 12'h5ac;
 filter_out_expected[824] <= 12'h8e0;
 filter_out_expected[825] <= 12'h655;
 filter_out_expected[826] <= 12'hb31;
 filter_out_expected[827] <= 12'h691;
 filter_out_expected[828] <= 12'ha4b;
 filter_out_expected[829] <= 12'ha25;
 filter_out_expected[830] <= 12'h74f;
 filter_out_expected[831] <= 12'hd18;
 filter_out_expected[832] <= 12'h71d;
 filter_out_expected[833] <= 12'hb12;
 filter_out_expected[834] <= 12'hb4f;
 filter_out_expected[835] <= 12'h743;
 filter_out_expected[836] <= 12'hcf4;
 filter_out_expected[837] <= 12'h73f;
 filter_out_expected[838] <= 12'h9e0;
 filter_out_expected[839] <= 12'ha33;
 filter_out_expected[840] <= 12'h6f5;
 filter_out_expected[841] <= 12'hb39;
 filter_out_expected[842] <= 12'h68a;
 filter_out_expected[843] <= 12'ha1f;
 filter_out_expected[844] <= 12'h752;
 filter_out_expected[845] <= 12'h967;
 filter_out_expected[846] <= 12'h62d;
 filter_out_expected[847] <= 12'h9b5;
 filter_out_expected[848] <= 12'h5f0;
 filter_out_expected[849] <= 12'h8f2;
 filter_out_expected[850] <= 12'h672;
 filter_out_expected[851] <= 12'h933;
 filter_out_expected[852] <= 12'h5a3;
 filter_out_expected[853] <= 12'h9cb;
 filter_out_expected[854] <= 12'h56f;
 filter_out_expected[855] <= 12'h8c8;
 filter_out_expected[856] <= 12'h6d4;
 filter_out_expected[857] <= 12'h6c7;
 filter_out_expected[858] <= 12'h88c;
 filter_out_expected[859] <= 12'h524;
 filter_out_expected[860] <= 12'h8a4;
 filter_out_expected[861] <= 12'h43d;
 filter_out_expected[862] <= 12'h893;
 filter_out_expected[863] <= 12'h47b;
 filter_out_expected[864] <= 12'h7ec;
 filter_out_expected[865] <= 12'h5f3;
 filter_out_expected[866] <= 12'h635;
 filter_out_expected[867] <= 12'h8f5;
 filter_out_expected[868] <= 12'h52f;
 filter_out_expected[869] <= 12'ha2e;
 filter_out_expected[870] <= 12'h753;
 filter_out_expected[871] <= 12'ha18;
 filter_out_expected[872] <= 12'h817;
 filter_out_expected[873] <= 12'hba1;
 filter_out_expected[874] <= 12'h77e;
 filter_out_expected[875] <= 12'hd58;
 filter_out_expected[876] <= 12'h712;
 filter_out_expected[877] <= 12'hcba;
 filter_out_expected[878] <= 12'h9d7;
 filter_out_expected[879] <= 12'h9d4;
 filter_out_expected[880] <= 12'h49c;
 filter_out_expected[881] <= 12'h94a;
 filter_out_expected[882] <= 12'h955;
 filter_out_expected[883] <= 12'hbaf;
 filter_out_expected[884] <= 12'h66b;
 filter_out_expected[885] <= 12'hb08;
 filter_out_expected[886] <= 12'h6a4;
 filter_out_expected[887] <= 12'h7d9;
 filter_out_expected[888] <= 12'h644;
 filter_out_expected[889] <= 12'h70c;
 filter_out_expected[890] <= 12'h257;
 filter_out_expected[891] <= 12'h838;
 filter_out_expected[892] <= 12'h002;
 filter_out_expected[893] <= 12'h58d;
 filter_out_expected[894] <= 12'h18b;
 filter_out_expected[895] <= 12'h0bb;
 filter_out_expected[896] <= 12'h2b0;
 filter_out_expected[897] <= 12'h00a;
 filter_out_expected[898] <= 12'hfb4;
 filter_out_expected[899] <= 12'h4ea;
 filter_out_expected[900] <= 12'hdfb;
 filter_out_expected[901] <= 12'h60c;
 filter_out_expected[902] <= 12'h29a;
 filter_out_expected[903] <= 12'h3e7;
 filter_out_expected[904] <= 12'h809;
 filter_out_expected[905] <= 12'h448;
 filter_out_expected[906] <= 12'h8fa;
 filter_out_expected[907] <= 12'h7a9;
 filter_out_expected[908] <= 12'hfd3;
 filter_out_expected[909] <= 12'h9db;
 filter_out_expected[910] <= 12'h7fe;
 filter_out_expected[911] <= 12'h983;
 filter_out_expected[912] <= 12'h7be;
 filter_out_expected[913] <= 12'ha30;
 filter_out_expected[914] <= 12'h688;
 filter_out_expected[915] <= 12'ha80;
 filter_out_expected[916] <= 12'h63e;
 filter_out_expected[917] <= 12'h994;
 filter_out_expected[918] <= 12'h771;
 filter_out_expected[919] <= 12'h942;
 filter_out_expected[920] <= 12'h62a;
 filter_out_expected[921] <= 12'hb1f;
 filter_out_expected[922] <= 12'h666;
 filter_out_expected[923] <= 12'ha36;
 filter_out_expected[924] <= 12'h9d0;
 filter_out_expected[925] <= 12'h6f8;
 filter_out_expected[926] <= 12'hcfd;
 filter_out_expected[927] <= 12'h68d;
 filter_out_expected[928] <= 12'hae8;
 filter_out_expected[929] <= 12'hb61;
 filter_out_expected[930] <= 12'h6b2;
 filter_out_expected[931] <= 12'hd7b;
 filter_out_expected[932] <= 12'h7ed;
 filter_out_expected[933] <= 12'ha0e;
 filter_out_expected[934] <= 12'hc25;
 filter_out_expected[935] <= 12'h7c7;
 filter_out_expected[936] <= 12'hbdb;
 filter_out_expected[937] <= 12'ha9f;
 filter_out_expected[938] <= 12'h7e8;
 filter_out_expected[939] <= 12'hd73;
 filter_out_expected[940] <= 12'h70b;
 filter_out_expected[941] <= 12'ha12;
 filter_out_expected[942] <= 12'ha54;
 filter_out_expected[943] <= 12'h6ef;
 filter_out_expected[944] <= 12'hb0a;
 filter_out_expected[945] <= 12'h668;
 filter_out_expected[946] <= 12'h974;
 filter_out_expected[947] <= 12'h634;
 filter_out_expected[948] <= 12'h965;
 filter_out_expected[949] <= 12'h576;
 filter_out_expected[950] <= 12'h8e7;
 filter_out_expected[951] <= 12'h65e;
 filter_out_expected[952] <= 12'h6e5;
 filter_out_expected[953] <= 12'h98e;
 filter_out_expected[954] <= 12'h465;
 filter_out_expected[955] <= 12'h56e;
 filter_out_expected[956] <= 12'h388;
 filter_out_expected[957] <= 12'hac6;
 filter_out_expected[958] <= 12'h4d5;
 filter_out_expected[959] <= 12'h86d;
 filter_out_expected[960] <= 12'h811;
 filter_out_expected[961] <= 12'h672;
 filter_out_expected[962] <= 12'h9cb;
 filter_out_expected[963] <= 12'h766;
 filter_out_expected[964] <= 12'h684;
 filter_out_expected[965] <= 12'hd12;
 filter_out_expected[966] <= 12'h3e7;
 filter_out_expected[967] <= 12'he9e;
 filter_out_expected[968] <= 12'h702;
 filter_out_expected[969] <= 12'ha94;
 filter_out_expected[970] <= 12'hc48;
 filter_out_expected[971] <= 12'h7d3;
 filter_out_expected[972] <= 12'hc28;
 filter_out_expected[973] <= 12'hac2;
 filter_out_expected[974] <= 12'h892;
 filter_out_expected[975] <= 12'hc5e;
 filter_out_expected[976] <= 12'h6de;
 filter_out_expected[977] <= 12'hab9;
 filter_out_expected[978] <= 12'h67c;
 filter_out_expected[979] <= 12'h8aa;
 filter_out_expected[980] <= 12'h4cd;
 filter_out_expected[981] <= 12'h704;
 filter_out_expected[982] <= 12'h42b;
 filter_out_expected[983] <= 12'h4af;
 filter_out_expected[984] <= 12'h492;
 filter_out_expected[985] <= 12'h40c;
 filter_out_expected[986] <= 12'h094;
 filter_out_expected[987] <= 12'h785;
 filter_out_expected[988] <= 12'h110;
 filter_out_expected[989] <= 12'h7bc;
 filter_out_expected[990] <= 12'h372;
 filter_out_expected[991] <= 12'h49e;
 filter_out_expected[992] <= 12'h7fd;
 filter_out_expected[993] <= 12'h2e4;
 filter_out_expected[994] <= 12'h963;
 filter_out_expected[995] <= 12'h566;
 filter_out_expected[996] <= 12'h6f7;
 filter_out_expected[997] <= 12'h89c;
 filter_out_expected[998] <= 12'he9c;
 filter_out_expected[999] <= 12'h7e4;

 end // Input & Output data
//************************************


  parameter MAX_ERROR_COUNT = 1000; //uint32


 // Signals
  reg  clk; // boolean
  reg  clk_enable; // boolean
  reg  reset; // boolean
  reg  signed [15:0] filter_in; // sfix16_En15
  wire signed [11:0] filter_out; // sfix12_En11

  reg  tb_enb; // boolean
  wire srcDone; // boolean
  wire snkDone; // boolean
  wire testFailure; // boolean
  reg  tbenb_dly; // boolean
  reg  rdEnb; // boolean
  wire filter_in_data_log_rdenb; // boolean
  reg  [9:0] filter_in_data_log_addr; // ufix10
  reg  filter_in_data_log_done; // boolean
  reg  filter_out_testFailure; // boolean
  integer filter_out_errCnt; // uint32
  wire delayLine_out; // boolean
  wire expected_ce_out; // boolean
  reg  int_delay_pipe [0:1] ; // boolean
  wire filter_out_rdenb; // boolean
  reg  [9:0] filter_out_addr; // ufix10
  reg  filter_out_done; // boolean
  wire signed [11:0] filter_out_ref; // sfix12_En11
  reg  check1_Done; // boolean

 // Module Instances
  firfilt u_firfilt
    (
    .clk(clk),
    .clk_enable(clk_enable),
    .reset(reset),
    .filter_in(filter_in),
    .filter_out(filter_out)
    );


 // Block Statements
  // -------------------------------------------------------------
  // Driving the test bench enable
  // -------------------------------------------------------------

  always @(reset, snkDone)
  begin
    if (reset == 1'b1)
      tb_enb <= 1'b0;
    else if (snkDone == 1'b0 )
      tb_enb <= 1'b1;
    else begin
    # (clk_period * 2);
      tb_enb <= 1'b0;
    end
  end

  always @(posedge clk or posedge reset) // completed_msg
  begin
    if (reset) begin 
       // Nothing to reset.
    end 
    else begin 
      if (snkDone == 1) begin
        if (testFailure == 0)
              $display("**************TEST COMPLETED (PASSED)**************");
        else
              $display("**************TEST COMPLETED (FAILED)**************");
      end
    end
  end // completed_msg;

  // -------------------------------------------------------------
  // System Clock (fast clock) and reset
  // -------------------------------------------------------------

  always  // clock generation
  begin // clk_gen
    clk <= 1'b1;
    # clk_high;
    clk <= 1'b0;
    # clk_low;
    if (snkDone == 1) begin
      clk <= 1'b1;
      # clk_high;
      clk <= 1'b0;
      # clk_low;
      $stop;
    end
  end  // clk_gen

  initial  // reset block
  begin // reset_gen
    reset <= 1'b1;
    # (clk_period * 2);
    @ (posedge clk);
    # (clk_hold);
    reset <= 1'b0;
  end  // reset_gen

  // -------------------------------------------------------------
  // Testbench clock enable
  // -------------------------------------------------------------

  always @ (posedge clk or posedge reset)
    begin: tb_enb_delay
      if (reset == 1'b1) begin
        tbenb_dly <= 1'b0;
      end
      else begin
        if (tb_enb == 1'b1) begin
          tbenb_dly <= tb_enb;
        end
      end
    end // tb_enb_delay

  always @(snkDone, tbenb_dly)
  begin
    if (snkDone == 0)
      rdEnb <= tbenb_dly;
    else
      rdEnb <= 0;
  end

  // -------------------------------------------------------------
  // Read the data and transmit it to the DUT
  // -------------------------------------------------------------

  always @(posedge clk or posedge reset)
  begin
    filter_in_data_log_task(clk,reset,
                            filter_in_data_log_rdenb,filter_in_data_log_addr,
                            filter_in_data_log_done);
  end

  assign filter_in_data_log_rdenb = rdEnb;

  always @ (filter_in_data_log_rdenb, filter_in_data_log_addr)
  begin // stimuli_filter_in_data_log_filter_in
    if (filter_in_data_log_rdenb == 1) begin
      filter_in <= # clk_hold filter_in_data_log_force[filter_in_data_log_addr];
    end
  end // stimuli_filter_in_data_log_filter_in

  // -------------------------------------------------------------
  // Create done signal for Input data
  // -------------------------------------------------------------

  assign srcDone = filter_in_data_log_done;


  always @( posedge clk or posedge reset)
    begin: ceout_delayLine
      if (reset == 1'b1) begin
        int_delay_pipe[0] <= 1'b0;
        int_delay_pipe[1] <= 1'b0;
      end
      else begin
        if (clk_enable == 1'b1) begin
        int_delay_pipe[0] <= rdEnb;
        int_delay_pipe[1] <= int_delay_pipe[0];
        end
      end
    end // ceout_delayLine

  assign delayLine_out = int_delay_pipe[1];

  assign expected_ce_out =  delayLine_out & clk_enable;

  // -------------------------------------------------------------
  //  Checker: Checking the data received from the DUT.
  // -------------------------------------------------------------

  always @(posedge clk or posedge reset)
  begin
    filter_out_task(clk,reset,
                    filter_out_rdenb,filter_out_addr,
                    filter_out_done);
  end

  assign filter_out_rdenb = expected_ce_out;

  assign filter_out_ref = filter_out_expected[filter_out_addr];


  always @ (posedge clk or posedge reset) // checker_filter_out
  begin
    if (reset == 1) begin
      filter_out_testFailure <= 0;
      filter_out_errCnt <= 0;
    end 
    else begin 
      if (filter_out_rdenb == 1 ) begin 
        if (filter_out !== filter_out_expected[filter_out_addr]) begin
           filter_out_errCnt <= filter_out_errCnt + 1;
           filter_out_testFailure <= 1;
               $display("ERROR in filter_out at time %t : Expected '%h' Actual '%h'", 
                    $time, filter_out_expected[filter_out_addr], filter_out);
           if (filter_out_errCnt >= MAX_ERROR_COUNT) 
             $display("Warning: Number of errors for filter_out have exceeded the maximum error limit");
        end

      end
    end
  end // checker_filter_out

  always @ (posedge clk or posedge reset) // checkDone_1
  begin
    if (reset == 1)
      check1_Done <= 0;
    else if ((check1_Done == 0) && (filter_out_done == 1) && (filter_out_rdenb == 1))
      check1_Done <= 1;
  end

  // -------------------------------------------------------------
  // Create done and test failure signal for output data
  // -------------------------------------------------------------

  assign snkDone = check1_Done;

  assign testFailure = filter_out_testFailure;

  // -------------------------------------------------------------
  // Global clock enable
  // -------------------------------------------------------------
  always @(snkDone, tbenb_dly)
  begin
    if (snkDone == 0)
      # clk_hold clk_enable <= tbenb_dly;
    else
      # clk_hold clk_enable <= 0;
  end

 // Assignment Statements



endmodule // firfilt_tb
